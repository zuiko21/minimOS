������������������󓻱�9��K� I99��������������w������������������������������99�����D���A��[������������s�������������������������������1��91�D�K�4da9���������������w������������������������������3����4I4��I@LII9��������������w?������������������������������?��;�L9D��@A����������������s3w����������������������������s���9{�DFK�@DDD99�����������w7�7�������������������������������񿻱dKII��DDDLK9?����������33sw�����������������������������D4�96D L999����������wsq7�����������������������������;���D��1��LFDLk���������������933s���������������������������1�;<FiI��DDi��9����������3w��������������������������1;[�9��aD��4��DF����?��������1133�������������������������3����4KIN���DlDF��������������;41s�������������������������I��4Li�F�i4���FDDD�??��������{1A33�������w�����������������C�3���C�DiIa�DL@F�����������73DI77��������������������������I?�K���IDaKcK;4`@DA1������������d3w������w������������������C���4Dd��IC�;D@ F����������36AA77������������������������1�I9�iDa�6���D@ @L���������sFC3������s����������������{�C�4FD��?��4@@FC����������q3D3s�������s3��������������?�9i4�iLDL93�?��D  DA����������A�Cww�����1��������w������AD4�dFDC;����dD�{��������FDd7�������sC������33�w��73�<�FD@6��@i��?���DDF�?�������wdD3���ww������;3?3?1��FD�aaD�;���6DdD����������4FD7������sa����;�1191;�39�DDFK@F???��d�@D?��������4Da1s�����3;1113�111�1?1��4l��d@A��;���3Dd@��?��������6D7������s4�91;;44��39;DDD3L@FK;�{��dKDDi���������tF3w������w1?�3�91CAi13�?��DD�9d@DC�;����;C@������3Da3�����s3��9;1�I411?3;dFDDdd�;?{1dK���������tDD17����w?��114A�131�D DDc�FLDK;3�������a�7�������w6FC;sw�����s17�916�dDAa�K�C��@Dd93DFD��;?��{ K?��������1DI����w4?�aD4dAA14?13�@DDDC�dDD;3�������@A�?������w4FC37����s4?��IcK<d�Dd4C�@@DddLddD3��?�3@����������DDs����w���4�aCAAda�D4a;�@dDC;d4D���?��?�`������s4�d7�������s4o�1aa4FDDdaCcD@@Dd91D4��;{����?3�K�?������sDFD3w���w��s���aadAFDd1dd@DdFCCdd4D{���{?�����;������sDDDC����s47��4�AdiDAFDaAa�1�@Dl4;�;D������?��C;�����3FDD?��wdG�114Al1ddAD�CD�a@F�;1�d{�;�����s�A�������tDdCw����sO�KC�CFAdaAaFK Dl3�11;;��;��{�1i�N4�s������4DDDa?����sDc�11449aDddFDDdD@DF���3��??�4k�3�C�w������4DDdD7�����DG�3�3CAC�DFDD�D FCÿ;33;3�3�{d���?16�w���wtdDDD���w�wsdC111�9444DDaDdFF DD;34<3��34C�;��@K7���w6DdFD3�����sDA;11a3�A44i@4D@FC1�sC;;{3�D;��?�4DC1����w31DDDDA�w�s��DC��13�4AdDFDC@LD@D��{��c93;�C�3�����C137�s�FDDw���?���FD193�;113��C@CDFC3�;91C��6C33�� A�;7�w3DFDDdD7�����DC��931;���3`D@dF1dd4??dDFD ?�� C�K{w1dDDdDDC������dI{;;��1�;3����F Da�4DDDD43��D`   ??�@;1k?73DdCDC@C�����C����{��3��9;s��D@DF4FF@  D���D  D��@����DDLD4A������0C���?��{�?���?� �6Da6FD ;�d@����`9;<dFCDCD7�������A�{����{���[����@ �F94FDD3��@Dd�������;�;DDACDD7������4��������;{{����   a3K1c;d@k�DK����0;;1D@DKA�3DG�������C���������������@ 3K1c�@ ��dC3�����49y1�1�D DD41�4C�����tD��������������`  1c�d    C��;;�?���3�D D�A;sD�������������������� ;3�d    ;���4c�{�����9993�D Dd�sD?�����D����������������` �@ @  DC����13����� �99FD DA4?4��7��?���������������� ;34@D Dda�����������@;�9��@ @DD��C���s��D7����������������  94 d349;?����������d��A���4DDi91�{D�3��D���������������� ��4D3K9;3�������?����9{�K�񹻻��?�4?��1�D�����������������  ;{4�33K�����??�����;�1����������������D���������������� 3��;4�4�{����?�������������������?��C��1{Da���������������� G����;3K?�s�{3���������;9?����������A����dD���������������� k?����4;������;;���������C��������??�d�t�DD����������������  C����1K�?;?���C37��������������������?��a�DF����������������@K???���{������C;;{���������?����������O��C�@D����������������0A;{�?���3�{���A3�������������������{����1DD�����������������C�����;�13?����F3;{���������?����������D��D@����������������� a�{?�;�D�?����C���������������������D�D�D@����������������� F3�;���D������Da3;��������������������0�DA@D����������������� D��;??;3C��{?��dF3������������������C�DFD �����������������@F3;{�6A�����{DDa;�����?������������_���@D@������������������D;9?;;{9N{;{;�c�F3��������������������4D������������������;33�{36C3�131�1DD?�������������������D94@@������������������{93�4L496;�dC?���������������������D @������������������dk��93�CdDdC3��4C���?�����������������ID@D ������������������13�13dcD DC�?;4@k?���������������������d @����������������������3;D6DFD;��67��?�������������������D@ @������������������;��3dFC�FDD7��4D��������������������dD@ @��������������������1kfDDC1�Df?3d7���������������������d@��������������������3�DddkaK1��C�4���������������������94  ���������������������6dDDCa433Do�63�{�������������������@@@�����������������������@FD�1d�s�{���������������������� D��������������������91cd@DDaadDDk���c���;��C���������{�����;4D9���������������������F@ FDD@ F�?�1K?�����;����������������������������������������;cDDDD DFC3���c��������9�������[�����9�������������������������ddDFd6fk1��?;?�?����9�����������������������������������������44ddcDiF3���;;4�;������������y��_9{�������������������������C�DacFfF19?��17������K��������9��۹9�;��������������������۳444iCADlc���3�K�K��K�4����������������{������������������������CCF4�d6�?��3I4���I1����������ӱ�����������������������������6FC1FDÿ��{64K����DK�����������������������������������������ad��d�;?������k�?�DĿ��s��������?���������������������<�������Fc3�?�??;�c@;O���9������������?�����9���������������I�����9��4dD33�s����CD��?�������?������󽻓ӟ������������������������9�4FC�;;??;44K�3?������3��������9{�911������������������������DD3;33��1dO�1�K��������������9�����������{��������������FFCC�1��3��@O��;�O�������?�������DD������������������{?��;4Dd�a3�3d ����3��;;����3�������DDDd4d����������������񗷻۳O�CFDCd443�@���[3O�7�?���?�������DadID�����������?���?�9�;����4dCD4�FCCD 	���?����������������D�Iaad��������{�����;��������� CFDdFDDD�d K�1�������?�����������6DD�������������������D��D�dD4FFFD@�1�?��{��������������C4d������������������;99��;FFD�DdDAd ��I��9���������������IaFDD�����������������������dCFDFDdd@ ��F���K�;�?������������4D�D�����{��?�����������y�DDdFD�DD@ A��A�?������������������DFDd����?�y�?;3���{�;����DDddd O�F��������������������4�DDy?������3�;��1���������dFFDD@  ;?�D7�1������������������dDd���9113AAdc���?;[����<44DDD @D����L�?���������������Di��93C�4ididDI��A����������FDdD@ D���4������������������4��kCD4FAF�C{{���;9����DDDDd@D@D	���D��?�3?�������������C���C�d44aCCK�?���1������D FFD@d �K��K�i����D�����������������6443CLC�4aa43ӿ�A������ DDD@D3�K�����9d������������������a3C3C13��?��������� dd@DDKD@K������F�����������������cC�3C44443�3�?�?����  DBDD�@ @I������d������������������16313a;CF6��3�?������� FDDDK3  DdO��;���4����������������63CC�a3CCA;�;q9���������@ DDFD�D �DO1��?��C������?���������Da9c3446CF6���D�������@ dDk�@ �D�������������3���������DD13c443c1aaaCC�y494������@ DFD��  K�D������������s;�������Dd3CC41FF��0���?��D� DK�@ �4d��;�9��?���3?��������DDDa�C31ad1daad3������4I��@�@dcDD O�K����{��3g�����������FDD64CcCCfafC�ӻ����@���@ D�D�@F@Oa���4�����?��?��������DFCFC6acAcCAda�9[�;�4 ����0 DdK�@ D;�;����������?��������DDDaaaa64daa;���D  ����� ěL4 d����?�9������;�������tD 66a�aFdFddF�����   ����4 @a�K C1��?�?������?��������@@�acFAFAFFDd3���;�  ������ ƙ�@ �<�������������?��������@ 6adF4daacFC�� I�����6 I9�D {����9������������������  4FF1acD4d4dCFa�dI�����7�4  �D C�����������������������   Cd41FCFFFFdi0I�;�����@K�1 ��@ c��;�������������������D 46c4cFFFD4dDc�C�d��4��`�3@C0@ O�����K�����������������4D Cad4CDaddFFD6A��6K�����@6@�K�d �����A=�;����������������6D6addfDdddFDC3�����D 9`�C0D ?[���I������������������16