���������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ��������������������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@