��fk;;��;;;;���������������������������������?������������������;fFc���;;c㳳�?���������������{����������������������������=?�N$lk;3���>66i;[}���������{׽�{ߵ�׵��y��}����[�_���_��[��[}����;fNc�������d�fc��?��?��{?��9��������?������;S�?���������������3�f&n9;������fbn3��������dFc��y�����?����׻{���������y�����4�$ak;=;i;>nfk�;�4ddFDD`DC11�;{?���?׷�y������?��[�?�;?36�ffn;;;�㳳�d�b&;;�34dFFDdBFD$dFFD9=���������{�?����������3�3��6`lf���;3c�6�fb�;;DFDddFd@F@DddFF;=������{7�{߷�������f�fflfbd;3��;>f��"a�dddF�Df�FBDFFAa;?�������{߷������{;�f6�BfnFn6��;Fk;3�dbfcFDFF��d�F@lDdd$ddkC�����߿󳷷��{�����;�Ӷf�f��FfF�㳳>C��6ffa�dflD6afFd4FFdlFLF�D61����?߽�[��[����;3���fd�Ff�F�93���n;6lnl;�4k4�4�CF�dFDfFdFFaC;������?�[����9fckB&�db6f�F��;kf6��ff3FFFF4F4C4k4FCdfd3aaN6�y���?��;۹{;;?��dnFb&Ffd��ff6;k;<f6Ff��dda�<FAf�d4FFD�cFL4�441���?������fc��C�ffnd">6FNK9;;fnnf�3FFFCC�AFCDdafF�D43CKC�c={���{�9;dfK;�c�6F""fnF�>nfc㱶��ffC�af�143DF4lc�NDdC�kC�161l3�����3��b&����6F�"""fBb>dff�;;;6f�l;FKAk���cidcF44cCdD6�96�k33�9�1��f"$;;3��B  &�&B3�d�ic���ff3dk3CdCc@CAd4ND6d6�d3c�a1��3�;�6fbnc��ö6d""&fFb�c�ffk;��df��d�1<49fdn�a6D9d>��;3�3;n3�6��B &i3k;;Nf "nnF6>Fd㴳;3�l3�1�KFfa�FLacfDd�FC131f3��1kfNfB""d�n���b"""Ffb��f�fc>��fc<ca�1�C4I4;FdfIAcFD3>9c9;3a;3�>f6f"&4�n9;>F &fF>4�fin1��<i31cFcD<d644dKDacfƖ6�c333��3�3fFNFbfcl4c��b""*nnb��Fdf�k;3cc��C�66CDl4Fd6NFddC�;393;�3���ff>Nd,l6fn>n ffF1ffF�f�����44�cK>FCdd�Daa�CC�6�3��3��;9;fNK��BfcanfcnB""&fFb�>nfd>;63443C6akDdFDcdfF4d6�3c�;1�1?3�3�Ff;`dnndl>fb &nf3�dlncc��ikK;C�FFFF�d�d�iddKCF3Ó93�3�;�;9;n���L&d6ffc�" ""FNbnfffcƻ;��43CF�FDDfFFFF>aC3;3?;�;�?;3�63��D Lf�lf�f`"""�fBflnF�c�;;C�4�afF�F�ddCFC4�cF��3���u���{[1έ�@FBfffda�B" $f�bdf$f>;��3C�C6�ddiadFF�<4�44�a43�;s���?󳳳;;=4FF�nff""dd$"Bnccc����4<4fkCFCfN463CC�aF�s���}{��H@BnfFfnFb"b"ffb &F���;;13CCd1d44kDdfKD9cd3ca;31�;{�����@D@`bddfl  "�nB" fckc�<6�C�c3Kk1FF4Cc�1�99c�;{3{������y��@`D�&d�nfbb"""ffb"  ln6�9a��4dF��3C6dF�d91�c393�����?����q�9D@ BB&&fNd" f�B "f�kk;CafF13�fF4d3c;�����?�{���{�=4HD`d&Bdnff" "&fb`"F�kk;c4<4d�dc13cdFK>133;???[{����������@D F�bdfFb""FBd` fK6�c�KfFFCf;F;fKcd�61;9������{�{��??�@@d�&bf,ff�"""fn&&lfK3�4d44�aa4;<13C1i;3�;=?�?���{������9DB Bbff�F"$bF``fkf�3knFCda�cC�3�6��k3��5��?����������4LBD@.bFBbf"""b&fBf�$dd�3�aaacCCC��3�1�16�3;�����?������{{�D@d "jf�df""FfdfBNcin3�d6�d�cC;C����;1?�7�{?��??�����4@BD bf$fff�""" $nBnD$fNf;nFFCF�6;3cc�k;;?���7���{}�����$Bb  b`d�&   "&&bnFdfa3�CC�4ac1�a;kk>133�s�׻��������??[9D""&nf$`""" &FF�lkKc>�6�dCƴ6;Ccc11���3�;���??{��{����d� B�"dff" ".f1��4cC�6�FFf4cC9c3�����33�s�?���������{7�{@@�""*fnnB""&FF�9cñ�3�f1iC�1>1�3C13��;7�3�7����������=�D"""fd�Fb`""B�f9;9;KCd�F4an9c19k;;;;393���=;�7�߿���{}��`B  $"fffF""&�f��󱳓;1nFF4F>ac9>;�c1��;{��?3��??{{�??3F`"""""dnn"CF99;���1fCF�a6����;3;�;93���y���{_������s��D�b" "�nnd`" "ffnf���;93����46�6641���;3�?;??{�{��{������;s�3d " "&Fff$��K�9?���;96FF�6����3�;;3�?��{���������?;���nbbb"ff�b"""Ffk6;��;[�����aaca3;1;91�3�������{��{��������{��6F    &�>FBfK4�����93�F4���;�3����9;;{?���??���������3�?fbb"$fff""&ƶ;;�[��;����d>33�3��??������?�?{���������>d   fna�  f;9������?���;f9i;3��;�����3�;��������3�3�{bF".Fffb"ñ���ӵ�[���۹<aC63�;9�;;??3�������CC�;;{�����k;��<&$"d��Bd���{�{��?��{��CKcó�3�1�3��������?3�Dd39����{�3{3��36d" &fcf`"k;[����{��?99y96493Ci1�9�;9;{s���;�C;;�?��{������;��9f"dnNF"$;�{���?�ۗ����f9;c��ó?;{;�s�[�3�FDD3?���s3;�y?3�` "f6<`&ó�����;�3��91cAi6�C1111�1�s�?��s�d@ 1�����?���4�bfKKfb;?[_��=��1aC�n63�;;6�NFCa�3�;{{�@ di4K3��s�{��f�N6�FB&a9�����{�D�kcDi994DFFd;;;1;����{4d`k�;����3��??;f�;nb������=���<DDAD6�3C3Cc�;;FD4;;s�{�3NDD<�����{�;c����;�B$c����[�;DDAdAFFK;;3�D F3���?���CBF;������f3?=�ӳ���;�`&�9?��9�lFDl1�6F���94  @a�1���{{�d<;��������6ff�;{?��;�4�fc����1�91DDDID1�d�33K@FF�F1����;c���׿{����ffffc;{{;���di�y{�;1�DDLCDC�FK3f@dDdca�;{��6cc��{�����ffffff;?1�?���c;�F��DDDCL�fF��4�FNB@C�KF;{�����{;?�����fbf&fff����99���??�fFFDDFDAIAA�1�93�3k4a�1�;C?����;3������{��ffbfnffc���{�;{{��_dd�BDDDFD<1a�1c�3�9;;;KcC>;���;��7�{����?�&.f&ffffk[[����??�&FF�DDAK3C��;�1�1���4;<1�������?�{�������ff&bffbfc���;s�;[��``@DDDLd�ñ�f�1�;;39��3�;�����;���=��ffb�fffff?�?��{���DFDD�3c943�3��;9�;�1=����{��?������&�bbf�n&ff�=��9?���` @@DDDad���f�3��;��;1��������;;���?2f&f&&fff�fc�;�y���{�� DDdDD;a��9�;;��?��;cK;{��}����?����&&&`bfffffk;񷿻���??@ @@@DDDA�;dc;a�?3�{;�3������{;;??����6"bb&&&fffff���;_?�{�� @ @D�D33�43�;3�����6�;��{��������{���&bBbbbbfff6??;���?���@ @DDñ��K6ù;?;���1�??�����s;??{�{0 &&&f&nf�f3��;����� @ `B@@@d;;k�a3����;ci3�����[�3������2&""bbfffff��?�?��; @ D dD#���C�6���;;;C�3����??������b"`bb"bbbfffc{{;��y{�  D D&&s�C�i?�{�3�9;���;3;���b&&"&&ffnff����y����@@`@  @Db$c�Kc�3����;k43�����;;;�?{�"f"bb.fb&fcf;?�;�}���  @D@@@`$"k3�d9?d;{{93��;9;?���?�3?���  &bB&&fbff�a�����{{@`@@ $&b"C9d3;�9;3��;a�1��?��3;;��?�"""&&b&f�fffff��?�?��$@f  &���k;c��9;1�;1�;{��{3�C9?��`   bb"b&f�ffcd?�ӹ{�[{@@@@b&"$1;6C���;;3�;1����=���{c����""""b`bf&&&�nk?;��;�� @@b```";�d;�3�C1�;9{3����;3;?� " "�&&bbfffff����9;3�@ D $"""K;;K;?~7�6ldFld6fd;?�=�����b""b&"b"f&ff&cc�;3㱳�@@@F b"&"#��c{�;�ffddd���{�{��V& "b &b&bfbfn93�l3kc�BD @@@""34��y3{>;Nff�;?���?��bb"&""b&f&bf�&&c��6��>cD$Dd�$B   "  k3�C9�;1�31�d6>;?������6&f  " "&".bf�fb&c91�F9cödNFDDNB�b""$""C9��c����3�����������f&""b f&&bf&f��6��>3kNCKkdaF  B   �6�?�K;c>999;;y�����`&f&"`""&"bb"ffb"fk3kkk;>�1��C��4b"" ""C����F3�91333�������&bf"b&f""ff&fc��4��>CkKl��9� "  #<;=�?4dk3���;?�����0ff&" f ""b` &bb"�k>;i��K3>d69;;`"" "B" 3a�����FK3�;��w����@ &&b`"" b"f""f�"&cfac�;;��fffFۓ�bB " "!�;=�?7�c391�3�����4"f�&" & " &b "bb&fkkkc�;6�``"d�3�1 "  ""93���d��>9�;��Bfbf "&"""f "&f""fff4�����&&$&A�3�b b"    c���;q��C9339?��4 "ff&b ` "&b&& &nff��;ckKb$&d;�9`" "b$?;��;��;��?� f&b"""" &""b"&fff;������ bbF�;�f ""B$" "�;3�;3f3�?[��@@ "fb    b "b "&"ffnfc��[�9;f$&�c���  "  ""a�;���9kfd  @"$b"bb`" b &ffff;���=��&&�f�;0"" " " &�3{1;;;?0 &  &b  "$"&" ""&bnbffc�y����BBddkn���"" " " $1��?����ffb   "" "" &  " "&ffbnf��?���bbFF4�2"$  " & "&C;3�93��i�`"  f  "" &"&"bffff&fc?����$$f��9��" `&  " ia;7�?�c3B  """&  "bb & &&&&bbff�?����bNFf;1� " """ f3�}?� `"   "f  "  b" &&�bbfff�o�����Ff�3��9�" """ `""A�;;;��""  b"""$""  ""bb&�&�f6c����?nFa�����b"    "  $fCC3s���   "B"b""$"` "  $&fbffffc��{��cf�;�{;�  " """ "&C9;�;{�"" " "` " "" "&bbbfbfffk�����d�;[��?�b$""  FNF6�;��6  " "" "&" " b""&&&fbn6k������C����{��` "$"B"" &1�=�;� "   "` "& ""B`bbbfff3�����3�;�{��_�b " """ ifF3�;��0" bb"" "  "  & ""&&f&fff���׿߹��{����[B " "  """F��;��2 " "&B " "" ` " """b&jbff�������ӻ�{�4"" """$4d6;�?�`" & k� "`"  "   b"Bd&&ff��������׷��[�=�$ " ""&�>�s��b" " ";4" """ $" """"bf&&o����������;��3�;b"$""&"!aa6;7��_b "C " $"   ""`f&fff�����������{��?�" b cc�i;{�B"`  """""" " " &&"bbbk����������{{��{ӶB`" """&D�3�;?��� ""   "  "B    ""b�&.?{�������{_��{���4" ""46�;��B$ &" b    "BB$""""f?��������?�����?�$" " b"&Kac3���� ""  b "" "" "F`b""Ff�������_���y{�{���� b " "C�9;3����B " """ "  NFFKC������������󱱿;��6 "&"dacC��?�� ""B   &&fF$f�3�=;���=�������{���??d&  " "Cd�;;���"   " "$$D�,fFDf�1���??��[����9{������ """"B $��3��???�� "b" $"  &Nf"$d�cac;3��������������?��;4"    "3KC;??6"      ""d FFk6D��;[�����������3;�9���@" ""d4<3;3���{�"B" ""nFd�ÖfCcc;;?y�����}�����;9?;;�" b"Ckca�y{���DDB@  `f`f�4;4FF��;?{�������{{3�ӱ��6 " b  n9;1�;9{?0 "  F fFBFFdcK4�dlcc3�������}���