""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""���""""""""""""""""""""""""""""""""""""""���""""""""""""""""""",�����""""""""""""""""""""""""""""""""",�̈���""""""""""""""""""Ȉ������""""""""""""""""""""""""""",��Ȉ����""""""""""""""""""ȇ��������"""""""""""""""""""""""��Ȉ�������""""""""""""""""",��3����������"""""""""""""""""��̈�����h��3��"""""""""""""""",�s31�����������"""""""""""",�̈���f���6(��38�""""""""""""""""ȇ333���6���������"""""",��Ȉ����f6���b��38�""""""""""""""",��36ffh��h���b������""��Ȉ����ch����b��36��"""""""""""""",�s36b����33���3b������̈���h���(�a2���(��3f��""""""""""""""ȇ33fb���16c���1(��f����f�1h���(�a2���(��33f(�""""""""""""""ȇ36f(���ff1���16(��a6��c�(���(�a2���(��36f(�""""""""""""",�s3fb����h�ah��16(��a��12�(���(�a���(��3fb���""""""""""""ȇ33f(����6h�c��16(��a2��a2�(���(�a18��(�3f(���""""""""""""ȇ36b����16h�f��16(��a2��a2�(���(�a38��(�6f(���""""""""""",�s3fb����f��f3��16(��a2��a2�h���(�a3��(�36b�����"""""""""",�36f(����f��&ch�16(��a2��a2�8���(�a33��(�33(�����""""""""""��36b�����6,���c<�16,��a2��a2���a3,�a61��,�c3,�����""""""""",�s3f)����16)���c6�16)��a2��a2���a3)�a2c9�)�&39������""""""""-�36b�����16)���c2�16)��a2��a2���13)�a2c�)��c1������""""""""��36-�����12����c2�16-��a2��a2�1m�3-�a2f=�-��&3�����""""""""��33������12����c2�16-��c2��c2�31m�3-�c2&3c-���c1�����""""""""-�31�������)���cb�16)��c2��c2�3a9�3)�c2&c3)���&3����"""""""",�c3������)���3)�16)��c2��c2�3&��)�c2"c3)����c1���"""""""""�c31������12���6,�16,��c2��c2�3&1�,�c2�f1,����&3��"""""""""",�31�����c���2(�16(��c2��c2�3&a�(�c2�&1(����3f(�"""""""""",�33�����c(�ab(�16(��c2��c2�3(a�(�c2�&a(����33f(�"""""""""""�c31������1(�"��16(�h&3��3b�3(c6�(�c2��c(����36b�""""""""""""Ȇ33�����12#"��16&1(�a8�(�3(c6�(�c2��f(���36(�"""""""""""",�331�����c!2(��131(�f1f(�3(&b�(�c2��&6(���33f(�"""""""""""""�c31����c1b(��113(�"ff"��3(&b�f�c2��&6(��33b�""""""""""""""�c33�����1"���33ff(��""���f(�h�hc2���6(��336(�"""""""""""""",�331����36"���6ff"(���̈��"��(�ff(c2���f(�33f(�"""""""""""""",�c336��c6(���b"�����""��Ȉ����""(c2���&(�33b��"""""""""""""""�c331h���f���������"""""",��Ȉ���("b������336b�"""""""""""""""",�336h�����������"""""""""""",�̈���"�����33f(�"""""""""""""""",�c3h����������"""""""""""""""""��̈������336f(�"""""""""""""""""�c6��������"""""""""""""""""""""""��Ȉ���fc6b�""""""""""""""""""Ȇh������""""""""""""""""""""""""""",��Ȉ�ff(�"""""""""""""""""",�����""""""""""""""""""""""""""""""""",�̈�(�"""""""""""""""""""���""""""""""""""""""""""""""""""""""""""���""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""