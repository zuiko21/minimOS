                                                                                                                                  ������������������������������������������������������         ��������������������������  ���������������������������        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �    �����    �������    �    �������    �����    �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �����    �������    �    �������    �����    �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �    �����    �    �������������    �    �����    �        �    �        �    �                �    �        �        �    �        �    �                �    �        �        �    �����    �    �����  ������    �    �����    �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        ���������     � ������    �    �����      ����������         ����������    �          �    �          ���������                   �    �          �    �          �                            �    � ������    �    �����     � �����                 �    �                      �    �                     �    �                      �    � � ��                 �    �                      �    �   �                  �    �                      �    � ����                 �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �    �����    �����    �    �                            �    �    ��������������    �    �                 ������������    �    � � � � ��    �    ����������������������������     �    � � � � ��    �     �����������������                      �� � � � �                                                  � � � � ��                                                  � � � � ��                                                  �� � � � �                                                  � � � � ��                                                  � � � � ��                                                  �� � � � �                                                  � � � � ��                            �����������     �    � � � � ��    �     �����������������������������    �    �� � � � �    �    �����������������           �    �    ��������������    �    �                            �    �    ��������������    �    �  ��                  �    �                      �    �                      �    �                      �    �  ��                  �    �                      �    �                      �    �                      �    � � ���                  �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �    �������������    �    �                            �    �    �                �    �                   ����������    �    �                �    ���������         ���������     �    �����  ������    �     ����������        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �    �����    �������    �    �������    �����    �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    ���     �������    �    �������    � ����    �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �����    �    �    �������������    �    �    ���        �       �    �    �                �    �    �           �       �    �    �                �    �    �           �����    �    �    �����  ������    �    �    ���        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �    ���������  ������    �    �����  ����������    �        �    �                    �    �                    �        �    �                    �    �                    �        �    �����������������    �    �����������������    �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �������������������������������������������������������         ������������������������������������������������������                                                                                                                                        �