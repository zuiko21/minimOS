       ����D�D�NNKDDDDDD@@@@NKKD��ND����䴴���ᱻ@              AKK�NDND�A䴠
 �@���������NNA��DNNA������@              NN�DND���K�A�DND��NNNDDDN��ND�KKN�NNKK@              ��D�DNDDD�D��K��D�D
 ��NDND�ND��D�D�N@              DKND��NNNK��KK��@@D@�@ND����NNKN����䱻@              �D�DN@�D�N��N@ �@�D�D�NND��DNNN�DNNK@              DNDD��DNNK����A� �@  � @ D��D䴾��KK�NKN@              N�N��D���A�ᴻ@N@ J   D@@@ND�D���ND��ND����@              DNND�DND�䴴��@�  @ NNN �KDNND���ND䴾KKKK@              �����NJDNKKK @@  �D@ @���D�KA�NAA䴴���              NNDD�D�D�ᴴ��J@ 
 �  NN�  NDNND�NKKN�KDN@              �N�N�D�DNKK�  @ @  �D@ @DND��NA��N���KK�K@              NDNDD������@ N    �D�  �NDND�K���ND��              A�D�@ND�D�NA� @
    ND�ND�ND�D�KDDND�ND��KK@              �DND��NN��@@      D����NNNND�NNDND�KD�KK@              DN�NDDD�D�N�   �     NN�����@��ND��N�NA��KKK@              ��NNJN@NNK��@D D    D�_����D�ND�ND�NKNA�N����              KND�DNND䴴      �N@  �K�����ND�KD������KANKK@              �DKD���N @    �D�N������@D�ND��NDAD��KK@              NN�NDD�ND��     @NK��_������N�NN�N��ND�N@              �DD�NN@�N 
   K��������D�NDD�KDNDDDA�ND�@              D�NNNDDND�  @  @   N����������D�NND�D����ND�N@              ND�D�ND�@  @@  �D����������NNND�D��DDND�N@              �NKNNDND�    � �NK�������D��A�ND�N�ND�KK@              NDD�D�JD䴻      @仿���������DND�ND�����A��              D�ND�ND�N�D D  N@  K�_������N���K�NDKD��@              �DDNDDDND�    @   ����������ND��ND�KNK�KKK@              D���JN����D   � DK[����D�����A�KKD䴴�@              ���NDDDND��  �@@�N�����N�NNNNKKND������              �KD��@�N@ 
N D�����������D���KNN�KAN@              D�D��D�D䱴  @ @  ��[�A�A��ND�KD䴴�N��KNK@              A�NDN@�D�� @� @  JD���D��K��D�ND�KD�NKK@              NNDD��DD�N   �  N�����������D����N��A����              �䴴DNJND@    @@  D�����������ND��N�D�K�D�KK@              DD��DD�   �@   �A�����������NDK���N�A�@              ��KDN�N@�@  @ ND�������D��NN�DA��NKK@              �KDD�DD� @ @ @ � DNDD��������O��KDK�KNN��KKA��@              KD����K@ J  @�D�D�������A������A����KKDD���@              NNNDNDN@    @@D�@DNDD᱿�������KD�KDD������K@              D�D��D�� 
 ����NA�����@���NA��K�KANNKKK@              �ND�JAN@     K@K@@K���������DKD�DN�D���䴴N@              NKN�ND�D�     @@DD������������N�K�NKNNN�@              ��N�NDD@  @ D    �D�D���������D����N��A�D�N@              KD�ND��   @ ��   JDDNỵ��������D��AD�D�DK@              D���@ @        JD����K���䴴��NNN�D�D�@              �ND D�N   @D@  D�DN�����������KKD��N��N@              D�A� @��@@  
    JD��������������D�NN@              N��DD�@�  D @ND���[����KA�NND�N@              �D�  �D�D@@� �DD@�JA����_��K�K��������NN@              N� @@@DN@N@D���� ��@DN������A���A�仱����D�D�@              �D   
NNDNDN���D������K�KK������DN@              N  J�D@@D���O���NDDDK�D����K��KKK������N��@              @� @@��@D����������D�N���������K�������D@                @ D�DD���N@����KDN@�@A�KKK�KD��������NN@               � ���NDND�A������DDN� DN���������[�@               @�@  @D @@DN�ND����������K�DN�������N@               � @@
JN@NDND�DOK����NO�@ J@K��N��������D�@                �@@@�D�NN����NK��O�D@J���ND��������NN@                @@@ �D�D�A��@���A��K� N�D�K�������D@               @  N �NNKD�K����K������KD䴱���������@              �@ @ �DNDD@JD�DD�N���N�@J@N�NK��������K@               @ @�@@@��DDD�@�D����_�������������               @   D �DNNN@@�D���������� DD䱻������D�N@               �
  �@DND�����ᱱ����� DN���������KD�@                @J  @��ND�@@D�@�KN��� � @N��[������NNKK@               @  
 D@DN�NN NNO�D�D��_�@�A_�������DKA�K@               @@    DDND�@ D�K��������@���������NKNNKN@               �
  DNDND� NNK���������@���������D��KD�@               @@   
J@@@@��NK D��������� ���������D�ND���               @    D���NDD���������KK�������D����@                @@  
@ ��N�N D��������K��������NNNNN@              
  @@JJJD�D@D�ND@NK������������������A��KKK@                @@  D��D�NN�K����������������N�NN��@              @    @@@@@DN@DD�D@NA��������D��������D��NAKK@               
D� 
���NND��K��D䵱���� ��������N��NKN�KK@              
D   �@@@@D�@NDND�D@D���[���NDK�����A䴴�N�@               @@ @ @@��ND�NN@JN���[�@ @N@K����NNKKN����               @��
@�@�D@��ND��������   @�����������N��@              @  @ @��@ND�KN K��_�� D �@�K����DNDKND�KKK@               �   @@�D@NDND�A����@NJ@N@������JDD��N@                 
 
@@JJNJD�NND ���� DD� D�A���DDJNDNDNK@               @   JDNDND����� ND�@�D�O�NND��D�����@               @    J@�@NDD�D@  ����  �D�@N�D��DD�NDNDN@              
@� @   @��@��NN� ��� �NNN@�NDNDNNND��KK@                  @  @NDDND�D  ����  D�DN@�NND�D�ANNNK                  
  � @@NDJD�NND O�� @ NNDDNN��NNKNDD�K@               �@ 
 @��DND�ND�N ��  ND@����D�NDND�D��NN@              
@
   @ D @��NDD� �@D�  NN@@DD�D�N�ND�DND�K@                @     D
D�DD
N�� � D D��NNJN�NAND�D�D�NK@               @J @    @DJ@N DDND N@@� DNDNDNDNNA�N�D�N�@               � @       N@N���@  DD�D ND�JD��NA����KKNN@                   � D@�NDD�  ND���ND�@ND���NKD�ND�K@                      @  @D��NN@@   �D�@D��@��KNDD�K������              �        � @DND� @ @�N@�DNDDD䴱���NNNK@              
 @@      
@DD@��   N NDNDNNNDDNDN����@               @           �
�@@D @@ DNN ��ND��N��D�DD�뱻@                        D �@�  � �@DND��NKKNNND��ND�KK@               @            �N@@N@@@N@DD�D�@NKD�����NND�@              
             @ @ � D� ��NDNNND����KNK�����K@                           D@ �@ @�@�N��DNKKN�A�KN��                          �� D� ND N@@�@D����䴴�K�KNKK��@                           @@N@@ D��@NND�DND��KK���N��                 @           @� D  D@DND�D�DNKK���N�����K@                             D� @�NN@�DND�D�A��A���@                            @ DJ D   NDD��ND������A�K�@                            @ � NDDNDD�NADDDD��A��KD�                              D@ N@ @N JDND��D�������NNNDANKK                                 �@ @��D���DNNKK�����������@                             @  @� D@�DDD��K��KDDD�����DN                               N  DD � �@���N@�K�����N������@                              D  J@N DDDNK�������������NNK@                             �  D J@NJN��NO�����������K��A��                             @  �@D�ND䴱�����������������                              @N���ND�NKK���������������                   @            
D �@ND���NK���NK��������                       @       JJ@@NNDNDD������DK������������               @@     @       @D �D��N���������������������                �  
 @    @         �DD�NKD�������������������               @       @         @@ @NDD����������������������                  
@     @  ��K����������������������       