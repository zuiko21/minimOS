                         DDA����?�����1�4� D                                         DKFD����6;;�;�9����> C@@                                       NL��i��i�7;[���1D�D@                                   @D 4DA��3����l1�{Q��d���                                  @�AD���K�413���4K[����A��                                  �ęl����K;K�3a;ϳK{�ݱ�@                                 ADCA��l3d$�6F�9��;�4K��                                d�DF�K96KNFn4�gq;1��3���                               @LI�9d9A7�4`FdFB�FC3��K��``                            � @4�;�A�Dg�4AFdID3A6�ada�{�4�D                            D  �	3A�1FFDAd`ddbD�3`FDc;��A6�                           @D D�K��C��DFCADF?D341�3�?�A��@                      D  @FD�CN�01�1`1�3D464fl;����9�� @                    F DD4�A�1�FDK�0FID114Fc�3K4a�3?�� A�                   @FDDFA@I�D�4 A6BDC34F�413D���O4                    DDDDda@fAD��@ fCfC�N�CKC6�;������DD                   D�DlD@@DD4DFa� ��A�1�16d4F�3���c�@d                 DdCFADDD@$ Ad4DFA@ `	0 FCy6fD`d��3�3�;�aD                 ddDA�D@D@  D�  ��d9;�43ACF����3��7�;d                FI���B FFd F@Ad &FB	��d@;�443cddksk��u���              CDAf@4F� `k �4IqBFD@kA�1Dc���?����?�@`           @Ķ�D�DD�FA�   `fK�FA<a,��;C66���7?����;�d�N          DAAĖDII`d   $`C@6�?�a;3;3�������?�KC�         @`CCDFFIA@    FLa� �F a4fFa�ks�5��37���������F         `DD`d�D��     Dd@Dd@@DDf�f3K9�7�����\��D        @ d�CNA@    dFD�@4�C@`N fDnd6dI43�3��7�3����i�@        DDL44�D6      `4�@DFFD4D 343FKk9��;��������3CKc    @ @d�4aD03`  DF DFFBddDdd �d�da3;3w��s�;�����    @ @D�aN�FF @@DDCD DFdDD`dda `Ad�K�39��;�7?���w���D    ` dD@D�F4`DL`�4B4DDDFDAFDfD #343��ӛ������???�O�@    @ C0$C�9?�dFC@Df@D dDdDDD�fdFdFDdA�cnc�1{��?�������@     @1N�1�?1�DF CDd@�DDDa4dAf6IFDFCy��a3d43K��;�{�?������     `FĴ9�DDF4$D@@ d4�C>�3�3C�6A�~o9;3C33��=s?3;�?�;��k     dCF����` ddf@DB FFFD�1��1�3��4���C�36�C�??3{�;������     Nd�;A�9FFD1D  !� DD�cKK;3?;;77�6;�3k�6a1�633{;7���=�     df�1c1FF94B �FFC������s��?{7��99�1��1;?������<�     C�D�3�DK�@  Dfdi3;�??w�?�?3�s3��c��3;1�1���;�����[�@   @DD�D�C1Fd�F   F DFD�c37�����{���>�;4��c�;333�??��sy    DF4f���ndD@ DB$4nI�;��s���?��{w33�3�Fg�_�?�;;���D�   DL4��D�;Ff  `CDD63���?����?3334�9�3����������q�O�   	D4CA34�?3FcD`D   d�d�k;��������3;��3_9��?����?O�   <G�D��3f<aDD  `   Fd3��w�������{s93c�9���3���?�?��=q	�  �A1��caI$  D@ dddD7{��{�������?;3�KLa���9�������?�O�@�A����64a�d@ dDFFF$4���7���������;c4�nkG�6q1�;;�?����?@@�CCda�ÜCFD@DD@d@`$3;��7��������7��cS4���c���������@ �DCC41d6`D4 dFD@dd3{��?7��������3��3n3o�󷻳�����B@  �D41K>��DBF  dD`d N3�s{��������w��31vf�6��;������siN  NDd��9�K@a@4  FDFD$a67?�{��w�����?;1�K�s��?�3������� LDa�9�4`d�BF`   BAK3�7��??�������s��33?�6����w������O  dFI�k� 4`df@@   1;�������������?;�34���;��l;�3����C?aa�i<9�FDCCD0`  Ck1�s�3�������?��31�6�;��1���?������@�D��3�dF4$FC   A1fk3�CKCKs{����;Bc�<���m�[3;�������?���d4��C�Dd4`Af	`0   a�33dn�4D�c�{�?�4$D�fK�;{3�7�������{s1ddD�F��fdNfNF�BCB@  C6f7;;��C4?��6CA;K113�?{1s;?7���;@IK����1��FdDdD �`    d436;���{��37���C;337336Gw;�?������{ F�I�6�Id��Ddd4� `  KK3c36�f��?{?7��w��D&F7�4��3��?�������d�DI��f��1�D14dd C1 F  33;6d@$Ds??����   �;�F��;7��������@�DcO�1��CICF@Da0@` 33�3d   ���w��3�E;3�3������������6K���A�f @3@`D dfn����L���?;;�{����o?ys����������`DCK1Ñ��adfF4DD@ c��?�k ��7;;��;3�C;�o�;���3������a��D���kD6DF@d�CdfFFD4�;7?��6��W;����;�?k��9���;�_����@��CCK��9n�DddBC�1FD@dC3����;����3���??{�7���q�;?�{��������� �1�>CAddCCd�DDd3;{{?w����w�sw��{{�w�?�fK�sc7�=;�;����D�N�����fI4@FCDdlD6d`DKC����?��?�s�;��w77���D9��4��6�����F���9d69DDDCdDdCDddak7������??7�����s���&��c3�����7���3O��1���F9CF1DDDdFDb@dFfD9;���?�������??;{�;�6Ad3k3��?W��?���;6C��1��6�DddC@DF DBI1�������ww�{��?�7��~4�k����������;���;��I46FFF@``  $f3�����w�����w��?��ss46Fa3���3��7����������9nI�ND4 D4@4d C9���������3���?�??�?6Fdf;�;�o;ӿ����CA<;��A�l`fD   `  $�3��������;�������s�F�CA�?q��;{�?۳�L3��I$I Dd6`$C`@@D��?����w��?����?��vF1<�����������d1�C��4CFCAFFF0F DFi;3�����??s�s����10K�;7�;����?������c��CAI4`3�@4@$DN@dDFFC6;?������;�?��?���6�4a;;7�?�������?�N�9q�CFd>FC��`D @adFDF�63�??;����s?���?wsFcCG3���{�������944ddD3CFFFDBDdd$fCKK3s����7�K��?��3 dcF;{???��y���˽��6��4�CFc` @�`$FC�dL1a;;�����;3;3��??� $A1�;w��?{����y��s�9<d4�FDD@�@` Bfc34�;s����;�w7���s� D$c1{��s�9�����������F6Df �@FFCd�f3����w;��77����@FF�c7��;�;�7���?��ϻ�K1�Difd`G@` A$`4a�C3��?3�������w��7{�`Dda�c�;3�?�������;�4�cCKDdFLd4D+033��w{�??���?��3 BFc1f;3s�;??��?�}������9K<D9C�fd�dC `F6k14;;��?����~f6;?� dKa�3;3����{?���A�C�1ndkD`F dFCDa� C�;cs���ffcfbf�{4Dc�3���{�����=A9K�43�A4�D1�DdBFDd dc�1��3sf$ffff3��Fa44�?�[�����A@ᵛ�64DfC�BD$FKC�FC3c���w63;�3���w{0Df<K3?{��w3�������FI7����d3d1�dBa�6DcFFdC3C�7?�s3����s?{�`Da49�3�w??������D���39�D5`Fa44D4F�FC4dfc6�33����3;s;c{�3 DCCDo31��?�������oDDI�;�;�fKdcC� fdCCaaAF4;3�{w��33k>;7� "D�fq6;;��3ۻ������icKA��1�dc6A1�@DFFKA3f1��??7�ss;{;���6 BKD�63w?;�9�������D�6d;�33�CC3F�idC6dfddn1f�;����?����w�0BDdC13��f17��?�1��1F�ę�?61td1d��d�F�f4fFfC1F3��;�??w���;�@ Kc�;��4��{��>��A�K31g<FDccF�6F$;CCDCcKfC3�ws{?�����pdF$c�F3�?7��9��@I�FCCF��Adcf3IF;c14dfÑf4633??s���{wbFDdF`c34?�;�;�s����� �4d41DFC6FDc4�a��46i�D66�1c3���?���7�DddfF�c73�3�����4� C�CCFFddDF�94ffaadafC603�311;{;���7w�FCBDd��;��6Gw����;f ;a�44d4c�FFfCFd4f3dfFf366��33;�?7ww`@DfdfK7?��3?w?��y�䔴3adfKF;Cc�fFFfFDA4�>N��;333�7;s{�0a``dFf���s�3����;;�nafdD�`1ad6c66104nA�63?;?333;3FfF dddFAk;3�?7�����sO��;��c6FCdCAa14��DcFa3�3s6�3�37;�3�d1dFDFDD4d�c9��;�{����?O�C;l3FdDdd4facF3K�4cF4fc�339�{;���;�d��k@FdadfF1�1����?�����O0d�c1fDFCk��d��4�C3�{�s�;7���Fd�dfCFFdFfa4�33���;{����1O��C6a�CddDA6cK�;AKô3;3;s;�����;F9�dddD9�d;�6�;�?�?�����D�0?C�����DfFa�36>46���;�379�7;�?7�|AA�cFD9Adc�A�3333{?�����1����aS3�nACKAfc�3;3;4�3�3s33;�7s�3�d1CNC�@dD�4c�3;3{������;� @F�A��D4d333�����c;;6���3���?3�Dd�FFdd6c�;��?1�?�_��t��K`F96F4DdfF3�;����3��3�;����{���s3�Ai�FCFfa13��7��1?������K�@d9I�Da�1;�;3�;�36�3c��;�����;�3;�n46D�4l�K�;;;3�s�����3� @�C�d46c;�;;���3���;��63;;s����3s��a1CC;3�3733;�����13� 4Cd�K16�;37�{7s�?;6��7�����;�?���s<;KCafa41133�y��44�s�{���1�0 l44DKC33;���s����;3��?3��?73�{;���3Ddfdda6k�;;��sc93y���;DC@CCF9��33��;��w�{���3�����{;s�3���AD��CFFFdfl�;��3C��{9G?>F 4d�4�6��7??��7��?;7�7����w�{���;3cfFD1f�fF;�����3���3k��  l6FN��Kk;;������s�;��7�����s������4�fd6ff33��k7;�3���3  ddI4��c33��������?��{�7�;��{�?3�?�?;{u;0F��C�;�;����66��k �D��K3;�s��?{���?w��k7�?����;�7s{??�Dd�c�ca3�>���{O3a��0�2�3;3�{?w{����3{�3k��s�7��?���s��>;y��6c433?F;3��3�9�@D4@�C�3�?{�?w�������{�?3��s���?�w;�;��c93Cad{��?k�_Db1Fa�   �33�s??�������s�s�#�{{s{�����������<>�FK;k;33@d4�   d �33��?�s?���������??�s7s;7��?����s�n;3�K�1����9FFCdB   @k�6�3���?�����??���s�7���������;19;��D3�;��K� n@D    @�;���??��������?;������;�?7����??3�c�?�C4k?1���qy@  t4D    �3377;��������7���;�wsw;�;���������f?���F3��3?�;�   �D   �33��{�s������{����9�C������?������c���f�a3;��3   6�  o1>�;s�7����������?w�y���s�7{??���?���?;k�����C��6�    d40  �c;�?;7w�����?����?�1�?�?�{����������3;��4;�k3�35� @ L  �C33;;���w�?��?����{��{?ӻ��w?�{s�?�����3�?�a{�11�O�D        �3n�󳿿????�����������{������?������w33��F�s�c��        󓳳��{{��{��?��?��?|��?������������s;������K73���@       4�377w�?{���?��?����w����;�����������;��;�;ac<;;L�D@      