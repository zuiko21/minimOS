   �����������û�K��;��������������������������;�;������@        @ @D`C�Dl99i>�����;���9?9;[yy9���9��K��l��          $ `���a����F��a���;���������������>;;����ᳳF��K`       ``��NHfD4�<dd�dlK�=;�;�{����9�{9;;��˛��<;�<<��鶖�@       ��F��Hk�4d�˛H��[��;�9�����;�����?;9��;KIkÛ96���         l �`NB���F���i��������y{�������;9���;k�ᱶ��i�Kii@       @ NLd�Ll6�9�;�F�ỶK���9=�����9�;�����;��9;�i9k�<����        � d�NNC��a�;lk;@�d���{{���;�;;�y��;��<�ƹ6�;9��@        @�`NFLha�ƶ�N�� �?��������;������>9�����9l�@        �   N�NkD F�<a�K0�(��{��?;�������9���;ı�9���ki`          �D>���a仳��� ` ?��۽;�����9�����9����>�K<nCƖ�         � L+�	id�4�DdLl` � ����;�{9�;���?<��K9���kD���NKN@        d @�i�F��fƄ@���  dNN���������������;��L>Nl<a        ` �@� @Ld㓔i>�9;� ��  N4D���D�����ӵ�;�;���4ld��F�@        d�f�L���NKl��D��> ?�` �ll<���?>K9���;����<<c���N4�d        @  �Dcô��<�K����=� 
FL`K@���<A�����<1����<>D`�N�F�       � � f��lNKkN��,6K�鶖  d��l$�����K��������lKƔlF�K�         @�Ldi;4�d�;F���$a�i  �L,d;9��Lk���;�����ƴ��,ld�        `D`�〴��NN���l�KcL�;���d�F�䓖;`K�������<9ld��FKKN@         ��Nl<<$�KC��K9����@	��A�lD�n�kLi����{=���NldN@���l          L`d  Nll<��ƻ��F��~F�C��L6��K��3��ƛ?�lD�lFDlF@       `@$@ � �(dND�LNDDFNFN�Nn@��F䴖Ndó@����D�l;��F�L<lFĤ�ƀ       ��N�NfNF��l;�d���<l�`iD�K���l�ƻ��i��<nFĳ���l��B�nBF@       F@@�LN@JD䳓���K�K���kBK��KF�i;�������lF���ƖD��JD�l,         �`d�F�NlK�k��;��>FKL��~lld����fK��F�,;4Dn�Ll$Nd�F           ��<d��䳓�;��i�����O���dƻ��;�i����ll���dl`F�`�B�         $(`�l`NL`dK9�d��i����`�Ļ��`�䱹��F��=>Ld��D>����`�d�l@       ���a�@$Bl��lF��K��`�nF�?�LlK��i�ᶓ��Fl���<4��B���        D�d�ihHlF�NNL��N��yND�����F�9���Ɣ�K�N�NN<<��<0�`N         �l�d�@��<k˳��;ÿ�����c�����Lk�>na�ld�N�kIk�����@       N�N<�d����3�9��y��F�����NFľ���Ļ��F�@d�Ĵ�lNNK�?�       �a�KNFδ6�KI�FK俻?��l;<���ilK�4�@d�N�F��D�Knû;���@        @�@NDa>�<kNa��iK���<6ƛ������kK�D��@�FdND�;��>9������            ,$�K�ô����󻿴�Ki����Nl<dilF���;˳�9��������?@       �� nl�<<;K;�������lK�����DF�N�FLl�m��L9������91��`       d`N�Kl�B���K鱻���K��l;����N���D��?� ��9�����;�9����;@       ��!F��D�F��C��㹿�����4����CNi�斻�4�;��;;���9����@      H`��B�k`�K�9;���k���K;����NiC���9����������;��9���       >l;�l;KF����?�����������lK�;����� ;��;9�;�;���?�@         �kL<n��K�;�D���K����������ó�����< ��󛳿�;���K��?�        L�Ɠ�ka�F�N�K��۳�do��td����;�H;;���{�����99��@      ��.�LllLL�NNk���������������L;��;����ỳ�??��?�9��;@       L`d��FD`d�ƹ���i�������lA���ӛ���� ����a���K�Ln�N@      ��I��˼k9���K�� 99���Dn���L������<@������<F�ñA�@       �`d�9l>��9k��O�4����Lhi����K��ӳ��ii1<>���LakN�`           L����9�D�F����K�d���K�����9� ����㻓�nk�Ó���         ��$`BLnI�NNL<����C�?��FI������{��� o�����䳱�������0       Nf���ƴ�F@A�;����F���dl�D����������˓����?����������       DĒ @$�l滱�;��<���D��k����������N4l9;������������`       nFL, N<�K��;O����K�����������99;���K�����;������{?�       @��,@J�id�KC���������K<�����;�i���9���������?�߿��`       �DF N>L��ƿ�;��>��<F�No��Kû;���������������������       L䄄N����Dl���K��d�kC�O���K���{���������������;��`       $`Nh,<>DNL���K{K��n��@����;������������������߿�@        @dl(F�Æ�����i��i;;Ľ� k����d������������������{����       
 �n<�NND�����󖹹?� �O���I�;������������{�{�����@         @�`dD��d�����d���;�;��<���9?�������������������@         (LD ���.F�LK�K�{�� K?�������d��������������������{����       d�n�lln��d�O���@�@��lA���`�<i{�������������������       (ND�FND�F�Ld���LC�`�?��
L<@�ƛ�����������������������       D �nfhKNKF�ƿ�@���;ƿ��@d,� �����������������������@         ND���dFļ<kli��ù9�߰��B@ ��@���������������������         �$`Lf��nN@	n���;����$� D�K ���������������������@       � �B ��lHC�dN9���i�����B �  �� �������������{��������         `Nll@  `�鿿�����?�����` (�@ ���������������}����@        (F   �ƾ9�����������    �@  �������������������{��       F@    ��ƿ����?���9���  � ��  ���������������������@       BH  , L>�������9;��������   F@  ?���������������������        hNDN����������K�������  �`  ���������������������@        ����9�����󓛳�9;����    @    ����������������{�ן`         D�����������������������  N  ����������������������       ����;۳����{���?��������   n�� ���������������������`      n�;���{������?���������   �;�� ����������������������      �N�������������������1��   K�` /��������������������`       9���������?�����?���������   K��� ���������������������?�      �;���??����������������   �����������������������`      ��?����������������������   �4�K����������������������@      �;�����=������{�������;�@   �������������������?���=?�      ������������������������   1������������������������0      �;������{����������������   �9�������������������������      ��;{��{������������������d   
��;����������������������`      �;I����?���������������   <9��9��������������������@      ĳۿ=����������9{;��A���d`   Û;9���������������������;�      �;������������O��������?��   >�������������������������@      ������?�������K���������N`  �;;�����������������߻��@      �������?�����k[��������   �9��9���������������������      ����������������I{���k3�0  Lii9����������������{����?      ��?�����������������������  �仓�����������������������      ����������������ē��;;D�  ��ù��������������������@      ��9=?�{�����������ni9�;����  䴴n99��������������������`      �9������?��������A�;��N�  FNK���������������������?�      �����9�{�������9���a�;��o�  ��>ù���������������������`      ������{�������<�LD�C�9d��  @NĻ����������������������      �?[�����������K�� �9�ƛ�  ��k�����������������������@      ����{���������4���� a�l?�  iNL������������������������`      �9��{��{����������� �ô�K����$a���������������������??�      ��;����������������@Lik;���lH�����������������������@      �9����������������`$�ñ�����d��999�������������ӟ�`      9�����{����{��������N˻�� � �99�������������?����;�      �;���߿����������;KlNli1ilF< �����I����������������`      ��;{?;����?�������;������� �� l�99���;���������}����      �;����=?����?���{>��K NIC�@@`,`����9����������������_�      ;���=������������@<>���C�L��N@�ii>����������߿��?��׻�`      ������������������NB�Ld��� �N�Kii9?������������������      ��;;���񿟷�����N<i9d����dNKB�Ld���ÿ�����������������`      �����?���;��{���������,fN<��  d����9���������{���@      <�;;���=�������lk<in ���N n@  KL1�;ÿ������������{��?�      �1���������?���6��  D�FNDd�L�   �d��K9;�����������?����@      ii�;9�������9���D  
F����Df   �N�ic�����?�����?�{�{���`      ��������?;�����4  ����L � �(dlNIk�?�����������?����      ��n��99y���=��   @��l`$    `F�����Û�������������ӻ0      �9a㓻�����9�      BD�   �@NfĹk�9�����������?�����      ��û�;��������      ��   BFd�kC����������[����?=9?@      ��9��99;;���   B ��  
  ����d��?�����������y�������`       <�c��鱻�����B    �d�  �BLl�kC�k��{���������;���      �4�9�K��;�h  �  � �  @D,F�6��������������?�����ӿ@      �nKkN���;��;�   � F�  L���;��˿������?���=9󿗻�@      lKKKi9999�;9��l  �@ � ��$$lD�óñ�;���?������������?�      �������듓������ $$ `` @$B�lKN�;����������?��y;�      �KK���k�9;��F@hH fh$LlNN4����������;��?�;������   