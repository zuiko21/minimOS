                        D@DDD��;��󳓓���D� D                                         DDD�a�9k9?9?;�y��� K @                                      Dd�A��Ó�aC����{��dDD@                                    D 4L�d�1��û;{F�o�;;�D���@                                  @FNDC�K�;944K;��=��I<D  @                              @DDD�L9��;;C�a4���;��D�@                                D�d�ñ����46�;M��S���l`                               DDƖ94C�4D�DidD;9;9���1���                                NNFK�D1FK�fDDdD1�aK1���A1DD                            @ @���94�D;�4ddK@�n@dF���;ôD                            D  �9d��ID�AdAddA��4dFD�=��D��                           @D Di�Dd6KC�FDF�CF;4D9a�C�}���I9F@                      D  dD�DÖA��a91`N��d�Cd�4A�7��}9KC� @                    D dD4DOl?DdN1�Di`>B9���@C�C���� @                    @D�D�F@O�aD��DA�@ ddA�C>F3K6af@����;0�                    DDDDdl@4�D0 4@ D�4�;a3�CIC���{A���DD                   DF�F�FDDFDDdd@N@ Fc�C�c���4CFD39?���4 �                 DL4�l@@@D aD4FD1` D@I4@DI?FKFF�C��3�4@                FDddddBD` � Da  dd4Di3��da3CCD49�9K��?�;D                DFD�d@ddD F@F� FFD�cDdK;D;FFDs��y3��6��D @            @�DD��@��I� @K KDK9D`@C1�ddC4�a�6�??������ D           @�d�4D44d  d 1`d;1Dc�d���F�1�3�;���[��CD�          DA��4�FD�@F    �DCA@A@K��a;49;�93�9?�������IND          `@lFD�FD4C@    Ddd�� KF a4FD�����K�?����?���D        @@ @ iDF4N@     FDC@�F�@@dFFD;;�3i<�;?�����D�D        Dd�D��Ka     DD49@D4aD@A 4FCCcCC6�������;�����K4@      @D��44d� @   F�4`ddD`F�F �4�d4i9;c�;�;��{?��4�İ     @ `�DFĐ`d@D0 FFDF�DdF@4@ C�C�FC911��{����3��1��    @DDDK�c4aF@@`dkD DdBFDFDdF@@cCF1a��3�;;{�1��?�����d    ` dd@F���NDDF@D4FFFFdFDFFDa$ @K99;�A;?�;�{�����=��k�     @ LFFI�?KDDF@�D �@dDdF@ddd�F�DD`D��a>�3�9���{���@    `CdD����FFK cDd@dFFDf�FF��D�4FfDk3��CKFa����������4a     DFD�㓓�1DDdCD@dId99;a;3C�c�k934�a������������;��     Dkd9���@FL``F@ ddF3CC6��9;��>c3��4;C�a�����3����A     FAF���9fD��d D` FKD<;1;;;{{�;3����;11�?;;�����?K;     IKiA9�FDFI4@ KDDL4;C��;�?�����;;1a�;;>�9c��?��3?����1K     CDF��F�   FFFdcK�?��?���s��;�1��1����������?9��O@   @�ld�d�óF�i4   A@dFD6�;;??�������{93963;99?;�9?���9    FDDI4C��Df  F`D4NA;3�����{{���31���;43���;�?������4�   DN4d4�����FD@  DC�d6����������{{{{�3;3�;13���?���O�   	F�D�Ôk�FDD`$   $FD93;;���������?3��?3���q;k��������   K4ak�i��A4CF  D   FdC;??���{������3�13c��1k������������  �A����A4>FD@ d` DDdDc���{?{��������;���4Ka�C����;��{�C� �dk<k�;D4K@F@ DDddd@i;??���������?�;1c�4��9;�;;������@ ��ÔC����dFD@FDDFD d3���?�����{����;4;?�;��������@ @�4FFK1KD11dd `FD@F�7�?��������??3�9;K1o�A��������FD  KD�9��I4dKD  Dd F;���?�������;3��a�����3��������D�  FD�a9DL4`$d  DFDda;;s��������?���a����?�4;?������� DFA�9i94��@cF@FN@   FDd��3������������??;�;;4?�1k�;���=����O dI49a�ᳱ4 DCDDF@d   a1;���{��������;1��?�91�1A?�������� �d<C�K�d<`fD6@ @ >3?3����{�������1�3F��;�;>��?����9� �d�1���dDdad�FD    C�c��;AD7����34Da�;d����?�3���;�4@�ICěCC�DK@cFCF@   d693Di66DdC3����1DDd34a6O��;����������DD9F����4fFD`0K@`   ;A�>C����;iC����6cC�K16�??;�?;?���9@�LA������I4dFd a`@  A6;?����3���;��1;�;�G����������@�A���D4�dDdF; d  �k3��c�3��{3���3�dDF�;�k�;�����?���D�@I�Yi9<�FF`K� F  �;4d@;;??{�;�@  �{6�;��?�����@�D��C��4dCD`Ba0D` d�;;;D  3�����00K;;�;?1���������l�d��;��@@i`D a�����Oa����;� �g�G�O�����������@DK1�KF�1�4dFF�FBBFf�;?{�< ��?{{{����C�{o�6;;�;��9?������CIFA��FdFF@CAidD`D3��7�9c�;������;3�����1;�9����?�;@��4��;�Ddd�FdDfDd�;??��;�3���;?����?��;9k?����;������ �k���CDDi4dF9d�Fdak;����?���;;�{{���3�F3��9;{�����?�@4���4�C�@FCDdFDdl` FF;??{��{s������3����CF;�÷�3�����3��C���i11ldF@FFdada@ddac�����?������{��{{�?�?4l1�c�493�3������1��q���KDdD�`FFDFFFF�c�{�����?;��{��;����C�;9���;��������d�}i13CF�DBCFBDdFBDd4�???��������?��?{���?�C3�{[?�;��;�O6������F�DddDdD$4 @B  C3;{������{�7���{?��1�FK9�?7��?���9oi9��AdF� f d4` d���������{{;s���{��{344d;���;��߱��CF��񱴱l;C@ Dd@ �F@;;{�����?3�?�?��?;FCC����3���{����L1a��A�DCF@FFF`C@ d BDl1;������;��������d9;�;s�?��???���d;9K4CDKA d9dD`d2 @`dF33�������7�����{��{3�Ca3�������������I��dd�FF4@f@FDFF Fdl<;7�?�����?����;{?d3dK9��;��1������i;3ӑFFFN96@D$@FF`dDFc3�{���1?�3��?{��@Kdg�;�3�������O��I1��Did1FDdc `adDFFlcKs���?�;;;?;{��� da4;;�?��������i4Ffi``dF@D d4$C9ac;������;;3{{��� CC�3����?�;���������dI6DF@�DF`BDfac6{{������??���?0 d������{;?�9���K��913�CF��dd`d @d`KFCÓf����{{��{?����{@dFD;3��3�;��������{K��FDadD d`D@FC0F1k;{?���{��{��??`Da1�?���?�����۱9431d�C�dFd�DdDf@FdC�1;c;;???����3?��� `C�;;1��?������?�;�ɴF4KDF1FCd`DKc;11������f;3fc;{� d;Aa�1�;?�?����I�A�43�k4d$i� FdfFF� CC�3;??�3f6ffBfc��FCd�1�;���??��;4aik�I�4@C�FDa96$`FB�4N941����d$dfCcf3�?2DCKK�;3?�������D@CI?����FFC�@@FAdFF4FFC;;3;?;6�3�3����@fac��;����?�����;�9��9�4F6diCdFDd�Cdidd43�6;{�;���3;?{@DN?{�?��������DK�i933Dl4Fi0fCc�FFCC;c3��33��33��� d6a;3;;񿷳�����;�D4C����Aa�dc�BdD4ad4633�;;3c;6;{� dd�N;��9??������Na�i93�3F6D��4`4cdFFFCdac���󷷿;��;��4 Dad�3;�{��?����FC���I;�ia�d;4kl6Dddda��61;;{???���B dFC6��3�C������1D�D��1�FDoFD6C��1dFFa�d3>3󷷷������d fDk43�34;3;�������CFa1��3DdC1��6DD;1�Cdad316F���?������F@dD K;47���1�?����`lddiD�DC4cDk�F�F`�4�FKd�aak7���{{��0DFBFFC�C����;����91� NAFd9FDda4c�3�Faaddd3a6>1;;????����� dddd`�d?93������ ��ND�4FC�dd�dD6�6Fa�CFFFF34k36aa;;{󷿷��FFDBFF����3�;;�����D ;1�FFDdF�6CdacddD;dacc�FC���;3�����?�@@dFdda3���;1�??����4C��DaDdAdi3�F9CCc64DFa�3c;3;3�33�?;;�0FDdFFK93��?�?�?��6�4D�DdifD�k;44FfaC3�93��;3�;3�41D dddBF@4c�91�c�{����O�D��FC�dDd3aci1dfCAa���;c�󳳷3�;4FFd0FFFda4����;3�?����[O��1��adcDdiD�C�;4dcCc�3�???;�3�d1�d`FDddd��;9;?�����O�A�D�KFDDFC6;;14443ac93��3��;{s3�FKDadfFFFDd36��;�{�������G��F��i�dfFdd��3>3�f9<;;3���??;󷻻sD�6Dd4aaF93����??{��;�L��A�;�FDFFd4�1�6633���;;;3���w7�CF�;FFNF��cCó���?�������@?��KD��4acdd3�;�63�i;;?6C�3�???��;d�ND9dDddDóa������?�����@K0A�a4aadDd�3�3�;;3��3��3?�;s���3w�dK1�fCD6c19�;�?����0�CC��CFBKk6�3�3�;9;�;s�33���?;�s�6C4�DFCDC;3�?91��9;�����d�d�C�a<d��;;;�;1�;6;3�14;{3��s??��I6�kCF3�i9�3��1i{������i� @i�F���33���{�3����;�k3�?3����;3�;IdkAida;63;�����;������� dK1aaa�C;��?7�?7��?���{�;3�;3?���A3Ca1kCF�1a��;y;4k9�{;A@@d�FDk�C�3�;{��?��?;�7���?7���?�����KKFDdad�39��?��9����NF��C�K�3;;;7�{��������{��{s�s3���CD4�44fdK3;y1;a9;;���1D`<Fi63�3���??��?;�77��{�����3334f�FK44ddC�1�c����O��  F4D����;3����w��?���;�������??{�󿿿��D4F�66k;3;�1��y6O�1  K��C4�3��s{{����?�{��;s?s��{���s3{{;;��a�Ii��4���<�L�K0 9D�Kqk9;3�?����������c�;{�?{��??��;?���Di;33a��C�;{�c�� �K��3�?3�{{�����{1;{�;{��{��s��;3?�F�;A��C{�?���a���1;`D@�cc�3�?���?����{��?;{?7�������;��1�c�4a�313���D09la�  ` �K3���??������{���󷳿;{������3��;ai3F?�;;?� �C4   �33�?;��?���������?��?;{s��������9c���������dfCdD   @OK93���{�����������?�����;??;�������13;;k4d;;;;�3�@C�    @��3�;��{�??�?{�����{;s���������?��d���K����;B  �>@    �3�;�;{{{�����������?��?;���{����{1c���ad1�;;?��D   ?9`   ��;3;??�������������;���?;���������;43��K3C�;0$  �FD  O�93���{�;{{��������1�;�����{���������9���3;k1c�1d@ @ FD�  �Cc;??;{�����????����?�{���?�������;3q��Lk>9��   d  �9;3;;?��?�����������?�?������{{��������;�?�c�3�;�O�D        �cC�����{���?����?�{��4���;���{?�?���{33��Di3�4��i�`       �;3�;????�{�?��?�������?�7�����{��?������{3�?�3K3����        ��c3�������{�����??{�{�3��{����������{�?�����;�D`      