qA11AqDq{{�S1q�����A1�Q;�3�����DDDS@D��;�DD�@D}1�41�{;�����131�{����4KQ���ۻۻ�{��1CDA��DD@E3��@@@ADD@3A1�Cq[{��{����[u�[�[��6D}5����������F��D@DDDDM��`@DqA��W�q���۵�[�;�[�W�[��}��������9�D�DD3KutDdD�F@Kt��;����������׵��AD11{��[����{���1�0DDD����DCDD;�DD;q{}1�����w���[�{����DqG����{��{�F�9L4D@�@9;D`��@DD��{{{W����uUD�����K�15�DCAADq[��ۻ��4IyD�d@DA��DD��@D�7����1{��W4DDA�1���{�AS��{tFDA5�q5����D`D@��KFDDAi7��DDs���w{C��q���A���UQK�[���1�TAF{Q{�WS� @� ADD�k�FDD;��K�dA;�}�qD���s[VC[���[�C�A4A�AA91D@@��DF�vѻDK���qDDE{�{DDA����11AA�����K�A@�dT94DDK�4�L�K��D��E�t{>DC�ױ���S�cA4{[����DqDC9@@�C�D��A���;D1C�@4A{Q��;���1�IQ��K�����9�4AD44D��K�א���[Dq��@DDA�@F�A1ۻ[�tQq4k�C��K�[���C�;��DaC�{A@�y0K��� @�1DG�19{����A1[�������[����1���4�D}��A {@DD    K411�1�����Cq1;�{��q��������������DFD  ��@   @  @KD�u1a{���qg�7����������[���	pA�I;��@@@  ���@ @  D4DFqq4�;QA5[���	pD�{����K����л���@D�1D@    �@@       dKKCWsA�3�4{���@DDD�K����[4��@AAD[�   D     �        DA�K{�11W�{��}uDE���QTD@DD@A��@@@          @       	<@K�{{51{qQD @DDE��DDD@D@@Q1@        @           C����ASDA1@dDD@D@[T @DD@@ @                  i3�;��AaC51�DAD 1D@DDD@A@ d@     @               A���9{{7�DDqDFDD@F @                           La���9;�������A14   Dd   @    C   =   1                 Di;3�91�;��׽�ۻ�u    D     @�  @@   D          @    D;;���93����{{�����S1   9   @ �@  @                  @ D4�����;3��۷����������D@                                   @��99{�{ۻ�{{����������                                    $ `FId�����}�{�����������׻t                        @       F  `c��{��ۻ{���������{���}���K����Ö�DdD    a�>       $��� FK1{�{{����ۻ�����������{{�{[{�{����;;;;;;;@;��      FC;;d�BF�CK�����������{������{���������}�{۷׷��[9;K{1�`   ����@ FBl;�ۻ�������{��{�����������s����۷���y{�������@   @D�i;;{d@CF;�{{���������������������{��������{{���w�[��;� `f�6k;=��FD>d��{�����{�����������������������{�������׷�{�>@  $�Fd�;{;{<��;����{���{���{������������{[�������{������S���B  @`B K;�����K4�׽�����������������{�������{�׻����}���w׻{�@   @��K;�{{@a�K�w����ۻ��{����{��{�������{�{�������{{��;��3��  ;�����{���K�{����������������������{�{��������{����׻{�[�`@  D�;{[���{0 fa�w{�����������������������{{�������{�{ۻ}��;�;@  �3���Fk��� �k=�������{����ۻ����������������q�{��{�{{������4  3�<;v�Ʒۻ�k6D37������������������{���{۷ۻ�;d;�����������;�  @ �3��{{{C�㓷��������������������������۳�k��{�{{{�{}��;0  �k�9�����;6FD��������{���{���������ۻ��{�;��;�������{��;5�@  d�f���;����F fK������������������������{��3{�����{��{���{�>@  ���;{��������FC{�������������������������۳{���������[{���   ;4��{{��{�{�  a�{������������������������;�s����{��{���{{;4    ���;��;{{���� F���{��������������������{{���{{������{۷�;q�    <;3���������@  d;��ۻ���{����������������CK{������{���{{{��6@   c;�;{�;����p   ����������{�{�����{��ۻ�C�{{������{�{����9�    �;a�;������  BF9{��������������{�����������{��{��������{3@   3����;{��0 dF�={�������������������������{�����{��׽�{���     ii�9>9��{� f�d;3����{��{����������}{�{�������{�{��{�{{��>@    F�@bƷ����@ FLn3�;�����{�����{������ۻ�{��{�������������{>$    �N;�������fD9;�{{�������{����۷��{{��{�������������}���d    klk;{���{0@if���ۻ{������������ۻ��ۻ����{�����������{�N@      Ó���{�`FDc;�����{������ۻ�������{������{��{�����[�D`       kf��{{�{� @�di7�{��{��{���{���������۷���������{���ӳ;<`        �;{��{�@ ``Fi{�[{��{��������{�{�ۻ�������������׷;1�F@         f��׷��`  ���{���{������������{����{��۷��{{y1�d@ @       L3;��� $ N3�{=�{��������������ۻ���{���{{{{���iF `        @ Lk3��@ @   dK{��}�׻�{��{�ۻ}���{��w������ۻ����LB@$        $ $d�;f`   d�[�����������������{�����{���W��kFD @  N `     l6�c��    dn{�����׻��������=�ӻ������{���@@@N �  `       FFDl``  � Nd;{׷����׻�������;��{��{}�{@ `   Ldd $ @`     l@BNdd   Fk<$KC������������������}�ۻ��;1�@FD� �$B@Dd     @  D`B   N   �7���������}����Fda;|;{��f4��BFdD      D   @    f    BFd=�������������iö��s��4FD@@D�F ` BN      h@    B    @   F㻻�{���������>3���4c6+{;9kLl``@ d      B        `   F�C������{������������滻����dBD�DN@` K@@    
@    $         `C$�{������{���;9{7���{��ld�d@`$@f         BNB@    d  `FFD㻻�{��������3�9;{���9dD@`$FDBD @        B�    @  $dfC׻��{��������<6��û���9d4d� @F@$$Nd$       @$`fD    d   F�FFk�{���������C��kK1��������@B�HdF@d@D    @  F �Df@ ` `  6Nda{��������ۻkia1�K{���DF @d&@dd$`      B@ d��   d $`l6FC���{�������D3��iC���s��` @� B�f��       `l` BFDf` j@ @ F FFD�{{��������<Na�c����Dd��dF�fDd`d`    `   @D$ dD�D`d`@l $in@cۻ�{�������d�C<I{���@  fbFD@   �    l`B nfFd> `@` F3f�ۻ�������C�d��c{���@ �@ FFFFF$`   B  0 �@NC<6ĳ�D @ `$N40�{ۻ�����4d�l4F�{��     lfnd$`  `  D    � d`&�l6N;�4`` @ c;fc����ۻ�����Dd�K{���4 @  DfCC�FF@`  $`@$` dFD9��;�{�F@`fFK3D��������ۓDlD{{{��n fF�2F�  @ � d DF$`;{ۻ��S��6 d��Fۻ��{{��{k;Dd�c����t�  Fdck3�FD ` 4 D $F�`�{����F ;`Ffd64$7׻{�����D���DN{���� �c��;fF@@$� dB  FdfFFk{���{��d k$�f��Fk����{}��KD@LlC�����  �f�c;3�$   4 N` &�d�;������ C�fkfFC���{����3��$D����� �Fa3���>D$  �FB@  I4k67ۻۻ�۶�B�Kka4`d=�{���@�&f�f{���{`f6��9;16`   � ldF c3F�{{{׻��4`@3D366��FADD@D 6F4�����la3;;s��@   `+� FF@�C�c;��������@`D&��F@f0    @DDK" n@F;{{���C��;s��>    A� dFl`6����������fC;46$K4D@DDDDD�b�`���{�3�;7��{F@  $ �  D6�c�{�{��}���6DdN6k`Fd;D@DDD�b& 7���{{�;{��0B   I=` D&F�a;�׻ۻ�}��d$kdF@ F;`DDDDDDLC$"@;{����k;���1;@ @@ N��$ L$f�n;{���[�����dFafd0���@DDDDDd��n`����{{3���s�d      A��D�B�FD����{�����vF$dk<`�3�tDDDDDDNDLc�{�{��9{y{�;@  F  99`d dD3Ff[��ۻw���{��Ddd3dfF;w�DDDDDD���F@g���{{3���3N@ @  C�<d �D;���{۷�{�{{B�3i`ak���4DDDDDl@�L �;{��{{{�s� �F   ls��ND`4dd�{{��{��۷۷ C�F4n3k7��DDDAD��K;@ i{������{�` @@ @  K�;v3BFL4d��{۵����w�`;>C�C���{DAAdD�L;�� C�{�{{{{�< �� @  3���`@$�FD;�}�����{���Dc4fFflk9w�DFD��{{@c7�{���{{ B�d@ `��1�`Ddk��������{�s����FLFF�;{4AA�D���s��{�{{���  �D,  C��9``fda`˷�{�S{{s�1�;s{� fdnc���DAa{��ױ03׷���� h J@L  ;�i6D@dk�k�[Ck���;;;3���6�$dNC��DCDD��;=��������@  @a�D�  �1���dC�Gd>3�3������7�{�6`d�{D۱K{=~ ;{{{�  j�@KI@@@����NdB@a��Ʊ�9;;1�7���{{��ddc�dDD��ķf� C���D�@ND�A � C�q9B�� F�4;;4có;;3��;{����{��;DA�ld6��N9 Ll�@� i� D@	;�4a���$K<C�;FN�;;1��;9{���{s��>�CID�Ald�;D Dl`DF�L``HA N@ ����}}6a�;9d�9���3��;3�������{��3DDdhNLdDD�$DI�H@d
B��@   	{c����FK��Fk1��ac�;;3����{{�������ACD���F��K4��K{�hN$,$A�    �9;���l;dk�6a����;14a7����{�{{4DDA{�yLd��� K{s�`D  @D�   @ ;���3;3��k��kK>;K3�;;fB㷻{{�����4�}��Lw��A��s���� @    �{{���9c�>F�kCF6�{3����D9{{{{{�{7�DD׻���K{{{7{{JL"�       ��=�{��3�9f�;<dn;94;{�����c={{s��4FC����N���÷<3sD�H    �    ;[���{��>FN3�F>1�ffỷs����F�;;;;;w���L{�G�{;~C{Ƿ��"  �      ��;ۻ�����4�d�FkDk4l ;{���FC��9s�;1{�={K�������378l �F       5;۵���������FN@�" "k����d33�;{d��@�[K{{w�C�3���@d�@f     ��{[{���y��i;0�4�$�����2Ci;3�33; ��1�Kq{;{t ���n`   ;�ۻ�}qDD8  D�D  D �N�{���`f�33��;DLD@ K{�D;w1@   `       ��={�� @       k� @@{�6�C3;7�CD 7{�� d    `d K=��DDD D@  @@�  G�D@ �D��`BFF���DD�;4 D@` @D @@   @ ��DIL�D @       @ �y, @ A�;� k7��;�1N>DId�     `@@d$@D@  ��I��@@��       FD @@  A��1dk>�;;A9kD���<<<   BFNNd�NF��FD@���D@L` @  �   F@ L D��K�1��;��;1I;dlld4d�Dd���A�Ĕ  @      @  lD @  a��9;;3�;�1��1�3� LldaiikF6��FL{D�IDD����        F $H@ k�9C��3������9�;@�F��93�9kDD�F�LA�l9�K4@       �HDL�FC�D���;;��;;6 Dd�ka��<4����F�DĔD���1��<@       @   @  �;�F�K9=3;����3���3�16�1aaFDJ@FD᱓�CD��@ FFd@,   D9;���9a�����{;9@$c�6��3�K<���d@�Ĕ�����DLDfC�Kn���3��c�㻳43}�;C�