                      DD�D @@@@ DDDDD@                                        NN����NK�NN@@뻻��N@                                    @  ����JD�D�D���D�   @                                   @@����@NK��������D@                                       A�K���ᱴ�KDK�O��D @                                    任��N��N��KK��KN@                                      ND��@KD�D���K�����@� �                                   @��N����K���ND���D� K�                                   @@D䱿�D��������DD �                                    �D DK��KN���ND���� @@K�                                   @@ @K���ự���D��N@                                     D���KNK����A��NK�� @ �                                  �� 䱿��ᱱ���DK�K�  @�                                  ���D�����������K�D� @   D                                  ��DNỻ��������A�� @@@@                                   ��@�N��A���������KK��                                       ��@@D������������N��  @D                                  ��� �������񻻻��D�N   @                                    ���D��������������� @@ K@                                  �� N���������������@  @��                                  ��� NK�������������D @ ��                                  ���D�O����������������D@ ��                                  ��K�@�������������@  @��                                  ��KD������������������@@@ ��                                  ������������������@  @��                                  ��N������������������D  ��                                  �D�������������������  ��                                  ����O�����������������D @ O��                                  ���仿�����������������N   ��                                  �DD�����������������D @ ��                                  ��N������������������N@ �                                  A�������������������D@  ���                                  �D�������������������@ O�                                  K�@����������������D�  K��                                  KD����������񱿿��D A�@                                  �@DK�����[��������D  K�@                                  �@N����������������  K@                                  K�@������[������D @@��                                  AD�D��������䱱��N@@ D��                                  ��D䱻�ỻ�������KKK��   K�                                  K@@��K������D����D K                                  K@������������䴻�@  ��                                  D@���������񱱻�KND� @��                                    DN�������KDKK@@ A�K                                   @���������KND��K��  N��                                  @ NK������K�NA�N@ �                                   @DNKDN��������ND�K�� �                                  � ND�������KA�DND�ND ��                                  D  @NK@N�����K��D��N@�@ K�                                  �@D�@DK�NKN�DN@DD� K�                                  NK��KN�NND���ᴴN @   D ��                                  �K@��D�@NKKNA�D@ D   ��                                  �@KN����DK�����  �@    @N�                                  ��@�����N@��K�@ N @  K��                                  A� KK��DD�A� N��@ @ A��                                  N�@ﱻ���D�K�@N�D    ���                                  � �@O�DDỴ���D �D��@@  ��                                  NN@��D   D�@��@@   @  ���                                  D N@O��  @ A�� �    @ �                                  ��@K��  ND���@ @ @    ���                                  @ D�O����  K��� N    ���                                  D� O����@�@���  K@ @   @D��                                   D@K��������� N��N�@@@ ��                                   � K�������������D��� D���                                  @@ ����������DNDN@@���                                  @@ K����������A�N���A� D���                                    @���������������A�D ���                                   K�����������K������ ��                                   N  K���������������D ���                                    K�����������N�����@���                                   D@ ����A������KO������ ���                                  � K����K�����NK����N@  ���                                  @@����������DK�����@@@K��                                  @K@ �����������������N@  K��                                   O� ����������������@ ��                                  @��������O���@������@  ��                                   ��@�������D���������� @ ��                                  ��D����������DD����N@ @��                                  ��������O����D�K���D@@  �                                  ���K����������N����N@ @�                                   ������������D����D    @K                                  ������������D��D @  �                                  O��D���K�����NDᱱ�� @ @�                                  ����N�����O���@@NK�ND    �                                  ���D�KD�����@ D��@@ @��                                  ���ND��@�����A�D �  �                                  �K�D��DD@����D �NN@@@@��                                  ��D�� ����@  D@DD   ���                                  �����@ ����  @   �N                                  �ᱴ�@@�����   @@@�@���                                  ���A��  A���@D@@   ND�@ O�K�                                  �������@��D  @KD �D�                                  KK��K���@��DJ@ K��N  �KD�                                  �ᱱ���������@D  ��D@K���                                  K�D�����@ANN  ��N@ �                                  N��뿿��� ��@ N��D�  �䴱                                  @�K������NN@@  ��KN@@O��                                  �NK���������@  DN���  O��                                  KK��K�����  ���D  K�                                  �D��A�������DDNNK��D @���                                  KD��KK�������NDDᴻD�  ��                                  D�D��N����������D  ���                                  NN��D᱿�����ND�D @ K�K                                  �D���KK��������A����    ��O                                  D���D��񱱻���NNDD @@@K�                                  �����N���A���@@   K�                                   ���� DK����KNKNN   @ ��                                  � � ND�����KKD@D @  @O�                                  �����@DN��������@  @  ��                                   K��@�������@@@@   @ ��                                  ��@A����DK�������� J@ � �                                  D@���D ������     D ��                                  ��� D�����D @ @@  ��                                   D��� NK������@@� @   ��                                    D�@DD������@@ @ @@ ��                                  @@Dᱻ�@@NN��D @     ��                                    ����@D�N��@    @@ ��                                   DK���� �NDDDNN@@@@   ��                                   @@�D��  D�D��@@    @��                                   DK��� DND@DD� @ @  @  ��                                   NNN��� NDN��D N  @@ ��                                   DN�� �DND�� @@D    @ ��                                  @@ND����@DNND�DD ��    @ ��                                   @�N���NDDDDN @@ @@  @  ��                                  �NK���@DNNNN@@� @  @@ ��                                    D����ND�D@@DD�  @   ��                                  D@@�N���ND��D�  @@ @   ��                                   �D�K����D�N @ @    @ D��                 