                                                                                                                                  ������������������������������������������������������         ��������������������������  ���������������������������        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �    �����    �������    �    �������    �����    �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �����    �������    �    �������    �����    �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �    �����    �    �������������    �    �����    �        �    �        �    �                �    �        �        �    �        �    �                �    �        �        �    �����    �    �����  ������    �    �����    �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        ���������     � ������    �    �����      ����������         ����������    �          �    �          ���������                   �    �          �    �          �                            �    � ������    �    �����     � �����                 �    �                      �    �                     �    �                      �    � � ��                 �    �                      �    �   �                  �    �                      �    � ����                 �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �    �����    �����    �    �                            �    �    ��������������    �    �                 ������������    �    � � � � ��    �    ����������������������������     �    � � � � ��    �     �����������������                      �� � � � �                                                  � � � � ��                                                  � � � � ��                                                  �� � � � �                                                  � � � � ��                                                  � � � � ��                                                  �� � � � �                                                  � � � � ��                            �����������     �    � � � � ��    �     �����������������������������    �    �� � � � �    �    �����������������           �    �    ��������������    �    �                            �    �    ��������������    �    �  ��                  �    �                      �    �                      �    �                      �    �  ��                  �    �                      �    �                      �    �                      �    � � ���                  �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �    �������������    �    �                            �    �    �                �    �                   ����������    �    �                �    ���������         ���������     �    �����  ������    �     ����������        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �    �����    �������    �    �������    �����    �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    ���     �������    �    �������    � ����    �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �����    �    �    �������������    �    �    ���        �       �    �    �                �    �    �           �       �    �    �                �    �    �           �����    �    �    �����  ������    �    �    ���        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �    ���������  ������    �    �����  ����������    �        �    �                    �    �                    �        �    �                    �    �                    �        �    �����������������    �    �����������������    �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �������������������������������������������������������         ������������������������������������������������������                                                                                                                                        