        UUP  PUU UUPUU         UUP UUPUU UUP                       P P        P             P   P      P                UU  P   UU   P        UU   P   PUU                        PP      UU              P UU      P                     P                     P                         UUP  P   UUP  P            UUP  PUUP P                                                                                                                                                                               UU UU  UU UU UU                                                     P  P                                                UU      P  P                                                  P   UUPUU                                                  P     P                                                  UU      P  P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            ww                                                              p                         wp                                   p                        ww                                  pp                        wwwp                                                          ww                                  wpp                        ww                                                                                                                                                              ww     ww                   p                                  p      p                 wp    wp                           p      p                 wwp    ww                           p    ww                 wwp    wwp                          p                        wwp    ww                          ww                         wp    wp                                                       p                                                                                                     ww                         ww                                   p                        ww                                   p                        wwwp                                wwp                        ww                                   p                         wp                                   p                                                                                                           