��DC���?1�44;@;1�CO;�1FDd1O;;?CDDd3Dd33�333313D314@40D@y?4i?�?�N��;@ �;1�����9�I?��O1�F�4dDO0I9�pI99;C��� �F@�����1�D[tC{CKO�a9�yF{���?a;FD$1�C�3�DdC�3A;d �d@D@��k�4C�<IG�C�d@C[1=�1���KlDk��FDdO3K� t�0F@??DC��{���KK3d 0 �4LDk�K�9��1��;;CdC���i;4dND�1c;N@�g@D ���m9���14CK<C� � a�O4G�K��?S�K?FF��i11C�DDd1�L1�a 4K0`N@??4�������7�4;�{D�4�;�3�;?���9{dD;�A�lda�A3�C�1�D���K?�;I��D�K4��;1���1��31�;���9�0�CCD��G��4NttD@1?�����1��L�0 cD1;󴷱k?�3???�s;׳���K�d4?4�DdF�D4	LO�O�?���OFK  ���A;{�1�19�;{��3��KKD������;FKdD�a�F@c41{�����KKDA���D�94K���41�ó?ӓs{1;C<CN�Dv;C DF�0Kf DD���K�?�34A��C91�����;3��491�7���۳�;;�kC��4�O�4D��DD4?����FL3L41D�ao9�;11�?3�;s�[���C�|D�3;�@C nL@Fó���;�D�3�@� 4@K�9�;���{y�7������;����4�q�DƖLdDDFD���y������I93�K@�d��O?3�7��C9?9{s����������;C�;|`A9F@D  d@����??��3C�A���4�4�7�����=;{?;���?;�9{��1���DDDd �N@�{�����3�Ks�KF7�1��?;?7=4��=���=�3�?��y�C�1A�4A@� DD@�������ֳA�C@�D��?��;;{?�;��{������1�C��Dl0D0 `C@19��??��;;�D�@41�?4�3�s�;ӓ�;�;3�s4G�A�F��K D�@@@�D@��1�����;;s��󳻳���ǳ=;��1�??��?����K;4K9DK9i��ID` D@N���{�����?����}[�;;?�;�����9}�?7�;{;��C�N4�43�FD� @@D@�����??;{;��;9���?����3�??19{����?�?�{7�3�<4��A� dFFD�y9;񿿱�;ӱ���y�9?g����9�����?�??;3�<0DDKK4DDA`C�Dח<{�y{ӱ9;193q��{{s�S�?11�_�?3���;D0�CD	1D�K 40��D�����������y�����93�;�߽����y�����?;�@D@dDC�dD�DL6D��1�O?=�O����������w�����;�����1�34�K����4�;4�L4ikAF�A�;��D;o����3�{{�{���?������{�{��;D�G���C���@D`C�CND�dD�L1��D�C��?�������??��?�������??����CI��1K0;@��DCKFDD?DD;0DDDdi��������?;��?����s����91�1@����3�@FD 0DKIFL�COh ����������{��=���{�?���;�??��1���O����`��d@�DFDDDo D DF���;?�����??3����������_��1?�9����D;�;D@�9DD@KCD D @D��s�����{���?����������;ӓ��;��;C�����`;s�F @DDaiCIiAD�@D dL�9�?9��?������{?��?��;;?�T�D@k��?{�;3L@�KD�	DDNDD C��C��C�������;�ӿ���{��O�3������c @���;�d��FKD@@`FABO�`N����9�����?���S��?���a���{��LFDO�{?�{6A@C41�`D@DD?�`D���4������;{������?4F�?{���a�cIG���dD�<N$K��;3�D@@K�`K?�9�?��?���?7�{���4d���9��0Do����@�ADg191�F� ���@�9�;������?��������K�6A����?�cDO�1�� F�4FLK91�1c�DN 91�D���;�;���������=���dDC�di9?�3���CKk��D;�Dd�C3D�Df  @{O�1��=�����{���?�?�K�������?�7NDG�O���4F�C399�aF�D�C1���?����?������������F�F�;�1��AKi�;3�doD`k3�1�D�f1������{�����?���������FD�A1�����C1CF������@6�49a4�k`KFK0@��;}��{{�����{�����?d`�ƛ���?��FI��?��6K?�d@�93<>A;4993Id{{������������?����?�d�d�i9?��?C�aC4�?󳴱�9DD3�9��d�k;F|@@��[������������?����?�tK{Ai1���A�i4�@��?�6�Fñ3��a;KC��C�D���������D�������1���1������C;Dc@??�3I{�D?;��KCCK4;<a�K@����?=���O�������?��{6������I� @ �?��;?4D���K1y4C�d���������D��������a��1��{��C�I4�@o����<i0C1�4aC���;� @�1OI�1K���D��������4���{���K?F�4@�?��3���C�@;44�la3{�KS  D@�O���9D �;;������9DD�[�a�Kt�K�����;4�;@D�4idA;��DD9KA�<�LD@Dd@@�{7�DDDd��O��O���{;D?����4�Dl1;?3�� DIIK��D�@ @ D����DD DA���4yI�3�{󖖳��;I����dDD���{D@@C�LD�� D @���0� �FA;�����;��1d?���II����FC;�c�D  LC��L4@@@  D@@@��4�@`	c������O�5������˛�d�CC�;��D @DDd�FD�D @D @@ �{�d@@@FA4�������=?���������i�KC�1K`D�D��Dd  $ @��?�@@�dN;��������������������ac�{<@@ @DDIldDD@@  @@@@@?��N@D DdIa��I����������9|�9�ĔAc���d4@Da�� @ @D  ��?CD�F�9�����K���������������Dd��3>�@ @D��DD  @  @ o�<@@@D`D��������A����I��DÙ��D1�Da @@@@D�DN  @ O�[�D@F��K����O�@I������D��K�NFCD�4�F@@DFF��D   @ ���KD D@D�������K�����������LD;CD1��@@DFD@@@ @ @�;��@@@d����ɹ����D�������˖�L4`DLd@FC@@Dd��Ld D    @ �{��0@@DF����9��� ���{������dLDDdD�DdD@@ @ ��<D�  lD����������@O�����[�I��4�`dD`DDD@D@@ @   @�9ILd@DNK����99�����9�����K���LD�@@FDDBDD��dd @   @ @��d�  @Da�����;ٹ��������������NFDD@F��D@L LFD        ���L@d9ۙ���9���F�������@�9��D��FDDD DD� �@@@@@  DD @ ٹID�  L�������O�D���������@��ɔL4�D@�$D�`@@l@D  KN  ��9FA DN���������d��������D��9d��iF@@ N  @�D@@ @94��  �����  F����9�D4D�����99�@����II�L@@dF  D  @DD@N @��  ���N@@�9���{�ۖ@ ���������D���F���D @@�D@ LD@ ;���@  ���4�@ ��������D A���������I@���I��Dd D @�@  L@@ �� @ ����a�D��������	�����������D��D����L@`D @@DD@FD I���;@  ����L@ 	�������D������������������D@@@B  @@  @ ��9;��@ ߓ�Dd9�O��������ۙ����Di�D�� ` @D@@ @F@F@ KA����� ����d���D��ٵ��ѹ����������`��9���D@DK  @ @K������D  ����O�DL�����������������ěI��C�@  @    D@N�ÖD���K @��FK�HF����ٹ�������i����@�<��˔D @@@  @DDƑ;IiI��9@�����DDDD���������ۛ������I��D����l@@@    @@@ @`D9K���KCANK@ ���D�`IKۗ����ٱ��9�鱛��	������D�@@@  D��4KiAD��� ����F�DDƝ��������ٹ�������9IND@` @   @�FKDCND�ND�N@ ����N@ I���۹�?����������	�ɴ��DD   @  D�dLCDLL�DDID O���A�d��ٹ�ٱ��������Ö��I����1L@D @@D�dD�lLFDLdDD�@@����ILdɽ���������������I��I����L�D�      DD�LA��lFDDD@l���9��@DD���9�9K������9ƛ�K������D� @ �FDDFDDDD D@`����iۙ��D�Ld��ۙ�����������ɛI������D @   ��F     ������9��@�D�����I��������<C�I������ I   @ NF@@D@@D @dND�����󙛛�d�I�������������������<�K�����D  D   @�Ld@�����=����L@KI������ɛ���������ı铙��<il@     DL@  �@F�@DdO���y�ۛ�KADL�߹���9���Y���<�I�������@L@@ @ @ @���O�?��K����{��������9������������KI���I<��D@  @@@��4�K�������ٻ���D@���������������Ô��K����IL@@   @D ��1�@O�9�D�O��?�9���FI������������������ɛ�����D� @ ��=�O��K���@������ϝ����99���I������NK�9���@@@ @  @@󓗹�4D1����C��?�{���ۛ�ә����������I�IA����9��D@@  @d ;1��@�价��������9����D���ٹӹ������<<�ᴹili����D@@�  @ C���@d��������ː	�������ۙ���������I���<�<Dd    F?�D KK9��;�� {��K��?�������������<��NI��������@@ @@  ��D  I99C;�=��;@��9���ϟ��������<���IK�K�����D@�   O�   C�K9����={��?3���@�ٽ��y�����9�������DI�����I`@D  DND  @  <��K�9����s�99���������ٙ��9��I4���N��9��D@F  @@       �C�9������9��Ĕ��ۙ��������əD���I�I�ɼ�����@D  @         KA9����D DK��N���������99��dLKÖI�����Ad�   @ @D�O����D    ��A����Y������������LDDLI����i���@D  @I  @  @ @@@��      ��˔����񙱙9��9�ᖙ��NDƓ˙����ilD  F   @@F� �      59�II�����������i�D� DI���I�D D  L  @@   DD D       g�DK������񙙓�����9鑔�<FD K�i����@@ a @   @ D@        K{4D@���ٹ��9�9����K�LD�������D  @  L @@@ @D         �D@  �������������������FL�I9���D @ �     D `   @   @  �34d   ����������˙��K��L<L	�������@ @               {9L   ۱陹���������D9I�K���@@  �       @ @@@  �F@   �휔��9�����������IDK������LL<d@@@           s1D  �O�������Ù�i��ÖNI����DDL@ �     @       O=d@ @ ����K������铙����4��D@�����LD@@  @   @      ��@    �I���������������<4�@���<` � �             s4@     �I��������iI��L4D˛�����@ @ 	9 @  @    7�@  @ D�ƙ��������9��ɖ�Ė���II�K�<�@  �              �4@  @ ˛������9����˙K�����iFFK���������@ �@ @  @ @  @  4  @ ���K����Þ�KI�II<��LDA��9�KDD  � @ @@         �@   O����I������ɜ�Ö�KIN���L����A��K�@ K