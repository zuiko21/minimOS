                   DDDDDA   DDDDDDD@                               DUUUUUUUUUUUUUUUU   UUUUUUUUUQ@                           DUUUUUUUUUUUUUUUUUUUT   EUUUUUUUUUQ                          UUUUUUUUUUUUUUUUUUUUUP   UUUUUUUUQ@    @                  UUUUUUUUUUUUUUUUUUUUUUU   UUUUUUUUU@    UUT                UUUUUUUUUUUUUUUUUUUUUUUU@  UUUUUUUU    AUUUU                UUUUUUUUUUUUUUUUUUUUUUUU   UUUUUUU    AUUU                 UUUUUUUUUUUUUUUUUUQQ   UUUUUUT    UUQ@    D@           EUUUUUUUDD                     DAQ   UU    DUUQ@          UUUUUUT                           @  UUQ@   DUUUUUQ          UUUUUUU@                             UU   DUUUUUUUU         UUUUUUUT                             @  DUUUUUUUUUUU         UUUUUUUU                               DUUUUUUUUUUUUUP        UUUUUUUUQ@                            EUUUUUUUUUUUUUUUQ        EUUUUUUUUUU                           EUUUUUUUUUUUUUUUU@       UUUUUUUUUUUQD                         UUUUUUUUUUUUUUUUP        UUUUUUUUUUUUQ@                       UUUUUUUUUUUUUUUUT        UUUUUUUUUUUUUU                      UUUUUUUUUUUUUUUUQ         UUUUUUUUUUUUUUQ@                   UUUUUUUUUUUUUUUUUQ         UUUUUUUUUUUUUUQ                   UUUUUUUUUUUUUUUUUT          UUUUUUUUUUUUUUUT                 EUUUUUUUUUUUUUUUUUUT           UUUUUUUUUUUUUU              UUUUUUUUUUUUUUUUUUU            UUUUUUUUUUUUUQ             DUUUUUUUUUUUUUUUUUUUU@              AUUUUUUUUUUUUU          DUUUUUUUUUUUUUUUUUUUUUQ                UUUUUUUUUUUT     DAUUUUUUUUUUUUUUUUUUUUUUUU                  AUUUUUUUUUUQ    EUUUUUUUUUUUUUUUUUUUUUUUUUUUQ                    EUUUUUUUUUU    UUUUUUUUUUUUUUUUUUUUUUUUUUUU                    UUUUUUUUUU    UUUUUUUUUUUUUUUUUUUUUUUUUUUQ     UDD@         EUUUUUUUUUU@  UUUUUUUUUUUUUUUUUUUUUUUUUUU@     EUUUUUUUUUUUUUUUUUUU   UUUUUUUUUUUUUUUUUUUUUUUUUU      UUUUUUUUUUUUUUUUUUUUUUUUUU   EUUUUUUUUUUUUUUUUUUUUUUUUUT       UUUUUUUUUUUUUUUUUUUUUUUUUUQ   UUUUUUUUUUUUUUUUUUUUUUUUQ       UUUUUUUUUUUUUUUUUUUUUUUUUUT   UUUUUUUUUUUUUUUUUUUUUUUUQ        UUUUUUUUUUUUUUUUUUUUUUUUUUP  UUUUUUUUUUUUUUUUUUUUUUUT         EUUUUUUUUUUUUUUUUUUUUUUUUUU@  UUUUUUUUUUUUUUUUUUUUUU          UUUUUUUUUUUUUUUUUUUUUUUUUQ   UUUUUUUUUUUUUUUUUUUUQ@      UUUUUUUUUUUUUUUUUUUUUUUUUU   EUUUUUUUUUUUUUUUUUUQ      APPUUUUUUUUUUUUUUUUUUUUUUUUUQ    UUUUUUUUUUUUUUUUQ@       @PEUUUUUUUUUUUUUUUUUUUUUUUUQ@    UUUUUUUUUUUUUUUD          @AAEUUUUUUUUUUUUUUUUUUUUUUU     UUUUUUUUUUUQD@            @@AUUUUUUUUUUUUUUUUUUUQ@      UUUUUQD@                    DDDDDADDDD         DDDD                        @ @