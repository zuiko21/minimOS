                                               """          """          """"         """"         "" ""        "" ""        "  ""         "  ""            ""            ""            ""            ""            ""            ""            ""            ""           ""           ""           """"         """"        """"""     """"""""""   """"""""""   """"""""""   """"""""""                                                                                                          UUP          UUUUP        UUUUU        UUUUUUP      UUUUUUU      UU UUU      UP  UUU       U   UUP           UUP           UUP           UUP          UUP          UUU          UUU          UUUU         UUUP         UUUU         UUUP         UUUU         UUUP         UUUU         UUUUUUUP     UUUUUUUP     UUUUUUUP     UUUUUUUP                                                                                                       �������      �������      �������      �������          ���          ���          ���          ����         �����        ������          ���           ���           ���          ���           ���           ���          ���          ���          ���          ���         ����      �������      ������       �����        ����                                                                                                              wwwww         wwwww        wwwww        wp ww        ww  ww        ww  ww       wp  ww       wp  ww       ww   ww       ww   ww      wp   ww      wp   ww      wwp   ww      wwwwwwwww     wwwwwwwww     wwwwwwww           ww            ww            ww            ww            ww            ww            ww            ww            ww                                                                                                         �������      �������      �������      ���           ��            �����         ������       �������      ��  ����     ��   ���           ��            ��            ���           ��           ��           ��           ���           ��           ��      �    ���      ��  ����     �������      �������       ������         ����                                                             �