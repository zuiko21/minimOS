f33                    wwp wp wp wwp  wp                   333330                       p p  p   p                     333f                    p      p  pp  p                       3333                    ww p   p pp  www                     3333                       p   p  pwwp                        3333                        p p  p p  p                      33330                   wwp  wp wp p p wp                   ff333                                                          333f"fff3333f33"ffff"fff3333f33"ffff"fff3333f33"ffff"fff3333f33"fffffff33333333ffffffff33333333ffffffff33333333ffffffff33333333ffffff""3ff333fff""fff""3ff333fff""fff""3ff333fff""fff""3ff333fff""ffi������������������������������o������������������������������ffi                        �    �o    �                        �ffi                        �    �o    �                        �f"i                        �    �/    �                        �"fi                        �    �o    �                        �f"i                        �    �/    �                        �ffi                        �    �o    �                        �ff)                        �    �o    �                        �ffi                        �    �o    �                        �ffi                        �    �o    �                        �ffi                        �    �o    �                        �ffi                        �    �o    �                        �"fi                        �    �o    �                        �f3i                        �    �?    �                        �339                        �    �?    �                        �339                        �    �?    �                        �339                        �    �?    �                        �339                        �    �?    �                        �339                        �    �?    �                        �3f9                        �    �o    �                        �f39                        �    �?    �                        �3f9                        �    �o    �                        �339                        �    �?    �                        �33i                        �    �?    �                        �339                        �    �?    �                        �339                        ������?�����                        �339                        �f33333333fk                        �339                        �"33ff333fb+                        �f39                        �f33333333fk                        �3f)                        �3"ffff"fff;                        �ffi                        �3ffffffff3;                        �ffi                        �ff""fff""3k                        �ffi                        �3ffffffff3;                        �ffi                        �fff"ffff"3;                        �ffi                        �3ffffffff3;                        �f"i                        �3fff""fff3;                        �"fi                        �3ffffffff3;                        �f"i                        �0      ff3;                        �ffi                        �       ff3;                        �ff)                        �       "ffk                        �ffi                        �       ff3;                        �ffi                        �       "f3k                        �ffi                        �       ff3;                        �ffi                        �       f"3;                        �"fi                        �0      ff3;                        �f3i                        �ff3    33"k                        �339                        �f33    33fk                        �339                        �"3f    fff+                        �339                        �f33w  33fk                        �339                        �"33   3ffk                        �339                        �f33   33fk                        �3f9                        �f33   33fk                        �f39                        �f33   33fk                        �3f9                        �f33  p33fk                        �339                        �f33wwwp33fk                        �33i                        �fff    f3"+                        �339                        �f33 wp33fk                        �339                        �f3f p  f3f+                        �339                        �f33   33fk                        �339                        �"33www 3ffk                        �f39                        �f33   33fk                        �3f)                        �3"f p  fff;                        �ffi                        �3ff wpff3;                        �ffi                        �ff"    ""3k                        �ffi                        �3ffw pff3;                        �ffi                        �fff  f"3;                        �ffi                        �3ff  ff3;                        �f"i                        �3ff pp ff3;                        �"fi                        �3ff pp ff3;                        �f"i                        �3ff   ff3;                        �ffi                        �3ff   ff3;                        �ff)                        �3""    "ffk                        �ffi                        �3ff wpff3;                        �ffi                        �3f" p  "f3k                        �ffi                        �3ff   ff3;                        �ffi                        �fffwww f"3;                        �"fi                        �3ff   ff3;                        �f3i                        �ff3 p  33"k                        �339                        �f33 wp33fk                        �339                        �"3f    fff+                        �339                        �f33w  33fk                        �339                        �"33   3ffk                        �339                        �f33   33fk                        �3f9                        �f33   33fk                        �f39                        �f33   33fk                        �3f9                        �f33  p33fk                        �339                        �f33wwwp33fk                        �33i                        �fff    f3"+                        �339                        �f33    33fk                        �339                        �f3f      +                        �339                        �f33       k                        �339                        �"33                               �f39                        �f33                               �3f)                        �3"f                               �ffi                        �3ff                               �ffi                        �3f"       ;                        �ffi                        �3ff      ;                        �ffi                        �3ff"ffff"3;                        �ffi                        �3ffffffff3;                        �f"i                        �3fff""fff3;                        �"fi                        �3ffffffff3;                        �f"i                        �3ffff"fff3;                        �ffi                        �3ffffffff3;                        �ff)                        �3""fff""ffk                        �ffi                        �3ffffffff3;                        �ffi�������������������������3f"ffff"f3k�������������������������fffff33333333ffffffff33333333ffffffff33333333ffffffff33333333fffffff"33ff333fff""fff"33ff333fff""fff"33ff333fff""fff"33ff333fff""ffff33333333ffffffff33333333ffffffff33333333ffffffff33333333ffff3f33"fff                                                f"fff3333333fff`             wp wpw p wpw   wwp            fff333333fff""                p p  p  p p                     f""3ff33333fff                p   p p      p                fff3333333fff"             w  pwww p pwww    ww              ff"33f33333fff             p  p   pppp         p             fff3333f333fff`               p  pw  p    p               fff333f3333ffff             wp  wp   wpwwwpwwp             ffff3333