""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""�����""""""""""""""""""""""""""""""")����""""""""""""""""""""""�������"")�����"")�������"""����"""")�����"��������"""""""""""""��������")�����"")�������"""����""""������"��������"""""""""""""���������)�����"")�������"")����""")������"��������"""""""""""""���������)�����"")�������"")����""")������"��������"""""""""""""���������)�����"")�������"")�����""�������"��������"""""""""""""���������������"")�������"")�����""�������"�������""""""""""""""���������������"")�������"")�����""�������"�������""""""""""""""���������������"")�������"")�����""�������"�������""""""""""""""�����)���������"")�������""������""�������"�������""""""""""""""�����"���������"""����"""""������"")�����"")����"""""""""""""""")����"��������""""����"""""������"")����""")����"""""""""""""""")����"��������""""����"""""�������""����""")����"""""""""""""""")����"���"����""""�������")�������""�����"")������"""""""""""""")����)���"����""""�������")�������"")����"")������"""""""""""""")��������"����""""������"")��)����""")���"")������"""""""""""""")�������""����""""������"")�")����""""���"")������"""""""""""""")�������""����""""����"""")�")����"""")���")����"""""""""""""""")������"""����""""����""""��""����"""")���")����"""""""""""""""")����"""""����""""����""""��")�����""")���")����"""""""""""""""")����"""""�������"�������"���������"""����")�������""""""""""""")����"""""�������"�������"���������"�����"")�������""""""""""""")����"""""�������"�������)��)������"�����"")������"""""""""""""")����"""""�������"�������)��)")����")����"")������"""""""""""""""""""""""""""""""""""""""""""""""""")���"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""����""""""""""""""""""""""""""""""�����""""""""""""""""""""""""���������������""����""")����""����������"""""""""""""""""""""")���������������""����""")����""�����������"""""""""""""""""""""����������������")����""")�����"������������""""""""""""""""""""����������������")����""")�����"������������""""""""""""""""""")����������������")�����"")������������������""""""""""""""""""")����������������")�����"")�������������������"""""""""""""""""")����������������")�����"")�������������������"""""""""""""""""")����������������")�����"")�������������������"""""""""""""""""")����������������"������"")��������"����������"""""""""""""""""""�����"""")���""""������"")��������")����"����"""""""""""""""""""�����"""")���""""������"""��������")����")���""""""""""""""""""")����"""")���""""�������""��������")����""���""""""""""""""""""")����"""")���""")�������""��������")����""���""""""""""""""""""""����"""")���""")�������""��������")����""���"""""""""""""""""""""����""")���""")��)����""��������")����""���""""""""""""""""""""")���""")���""")�")����""���)����")����""���""""""""""""""""""""""���""")���""")�")����""���"����")����""���""""""""""""""""""""""���""")���"""��""����""���""���")����")���""""""""""""""""""""""���""")���"""��")�����"���"")��")����"���"""""""""""""""""""""")���""")���"""���������"���"""��")����)���"""""""""""""""""""")�����""")���"""���������"���""")�")��������"""""""""""""""""""")�����""")���"")��)������"���""""�")�������""""""""""""""""""""""����"""")���"")��)")����"���"""")")������"""""""""""""""""""""""���""""""""""""""""""""""""""""""""�����""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""�����""""""""""""""""""""""""""""""""""""""""""""""""""""""""""��������")�����"")���"""""""""""""""""""""""""""""""""""""""""""��������""������")��""""""""""""""""""""""""""""""""""""""""""""���������"������"���""""""""""""""""""""""""""""""""""""""""""""���������")�����"���""""""""""""""""""""""""""""""""""""""""""""����������"�����"���""""""""""""""""""""""""""""""""""""""""""""����������"�����)��"""""""""""""""""""""""""""""""""""""""""""""����������")����)��"""""""""""""""""""""""""""""""""""""""""""""����������")�������"""""""""""""""""""""""""""""""""""""""""""""�����"����""������"""""""""""""""""""""""""""""""""""""""""""""")����")���""������"""""""""""""""""""""""""""""""""""""""""""""")����")��""")�����"""""""""""""""""""""""""""""""""""""""""""""")����"���""")�����"""""""""""""""""""""""""""""""""""""""""""""")��������""")�����"""""""""""""""""""""""""""""""""""""""""""""")�������"""")�����"""""""""""""""""""""""""""""""""""""""""""""")�������"""")�����"""""""""""""""""""""""""""""""""""""""""""""")�������"""""�����"""""""""""""""""""""""""""""""""""""""""""""")����)���""""����""""""""""""""""""""""""""""""""""""""""""""""")����"���""""����""""""""""""""""""""""""""""""""""""""""""""""")����"���""""����""""""""""""""""""""""""""""""""""""""""""""""")����)���""""����""""""""""""""""""""""""""""""""""""""""""""""")�������"""""����""""""""""""""""""""""""""""""""""""""""""""""")�������"""""����""""""""""""""""""""""""""""""""""""""""""""""")�������"""""����"""""""""""""""""""""""""""""""""""""""""""""""")����""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""