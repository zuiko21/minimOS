����������������������������DK��������;ND�������������������������������������������������α�[���{��{��4�C����������������������������������������������IFC����?����;�KĿ���������������������������������������������F<?�����������O��������������������������������������������N�KK;�?��������������������������������������������������������A`�K���ӓ����?����i���������������������������������������������F����������D��?�������������������������������������������@D9���������=���KKK�������������������������������������������D�N�K;�[���;=��9<<Cß������������������������������������������� ai9���������?���D��������������������������������������������@˔�{���[���9�;�9�;�����������������������������������������DdNak����������3�1�d������������������������������������������NL�K�����������;��K�����������������������������������������D�dK������������?�iaK������������������������������������������lL<9�������{���?�;�ÛD����������������������������������������LDd��=�������߿{���<4�K�����������������������������������������F��K9�񷛿���{���������?�����������������������������������������K�;��{?�����=?�;��K����������������������������������������D�li3���{���?���?���;C�����������������������������������������DDD���y���;����??����4���������������������������������������D,l㱳���{������s��û��������������������������������������LF�D��������{�{������3�<���������������������������������������d��KK�O1;?���?������;?������������������������������������F@K<��C�;;��??��{��;�;1;��������������������������������������DF�a��k��??��{�������K�;?������������������������������������4�	l;;4����;����������??������������������������������������0�@DF���kk9;������?���9�o?������������������������������������d@�d���;;;;���;{�{���=���a�����������������������������������@  @�a9k;;�{{������9��������������������������������������@@FK4�>93�?���?9?��;��O��3�����������������������������������`�L4�KC���{���;������?;���������������������������������������DCklfl;;�����;����?�����7�?����������������������������������$d�ACLFi;{?{��?�;���;�;���;6�����������������������������������D �4��Lc�����{;{�{;?�����������������������������������������F@LkNCNc�a�;����������?������������������������������������`�f�4���>1�{{{;{���;������?3�����������������������������������LdKa�Fó��?��������>1�����������������������������������������F@d�NKa�;;4����??���;a�?����3�����������������������������������lD��CKa�����������{�������������������������������������������Dlalll�����᳿;�����;>�?����{�����������������������������������Dk�fF?;;>;��?�������{�������������������������������������9<@��9KDlK�������?���;�?�����?����������������������������������dd4�d @d3��;?;?����3�|?��������������������������������������Nnk@  K����������;��{����?����������������������������������DFD��Kk@���?{??��;;���?����������������������������������<dlk?;>�o�����{�{;;;;{�{��?����������������������������������nF;���>FNC�a��{�����÷���;������������������������������������Fó������;�;?�����;�3�����;���������������������������������1ni3���9;?�ó���?���1�;�?���?=����������������������������������f��??�;��f�;���KCn�;����;?�����������������������������������f�<3��;����F����c�;��{���?���������������������������������Kiak9�������k?�;㻷���k�����?���������������������������������a���{�;����K���;;����������3��������������������������������� �c�;?��?��3������?;?��󻳿�������������������������������� @1�;?��3����?�������������3���������������������������������  �43��{��?;�����;a��?;??���;f�������������������������������   3û;�������;���K` ;������s�l�������������������������������   Kl3�����3�;;?��4�NN3�������3c������������������������������@   �ci;{?��������D��������o������������������������������    �K;������;����d�i?����{6o�����������������������������@    k6������93���������k����������������������������������     L4CK;;����?����������{���6������������������������������    fn���??0C����������;�����������������������������������@@   ��C�����l;��������������{������������������������������     fKl>;���toF����������������;�����������������������������D @  N4�4�;�󶻴;���������������������������������������������  B   FF�KN;�?;����?��������;�������������������������������� @L @  KD>f����;C;�����������3���������������������������������@ FB@   �.CC㳳�n�9?���������������������������������������0 F    3Clk;;;9;4;>���������;3�������������������������������@ Dd`    D�;;û��Ó;?����������{����?������������������������ ��@  3N3û<6�1�Nc���{;���{��������������������������������� dd    adi;;6��<d9��?�?�����f�������?������������������������dC�@   CKN6���N�a��û���;����?k;3�����0O�����������������������F�@ H@ �ca�;?�dc�k4c;{��������D������������������������������FCF@    3�F6����>�li?�{{c������6;?��@  ����������������������dn@@` @43�û��Fc��Kk;��;�����@�;��@ @����������������������DKDa�   FF<3��l���㓱1�c�����@c�;�@D @ O���������������������K49�;�  f3lf;�3�`kik���{K;���dKk���N@@���������������������d;�3��  AKF9���4�D;;k1���k;���; f3� lD� ���������������������9�6NF;@@ó1df;�9;f㱳����???���@ �i�@ ����������������������l b � cFC�ó�NdF�;?���c���� d�  D˴ ���������������������nbNfF K �`f�;dn$3������3���>F�0  F@   ���������������������`db,.B ;f@�������nd���{;����F� �D� ��������������������nj$fd  @�C�f?;9;K;�����{>3���0@F   FIn��;���������������������Fdn`�`B3c10Kk3�;;3�lk;{1᳿?;�n   ����������������������������b�hn 14�0d;1������df9�F9;;�`D  � K��������������������������fb�F&`B;31l�kc1��;?�i�NFó�9`  $��w�����������������������dbnbb@3CC0<a��??�;;;{�N;93�   ���������������������������lnkf�Ơ3��4c�;c��;����;1k;��@D   ���������������������������fc1�;f�43��F���;?����������> �  ?{�����������������������9;1�;`1344 fic��������{;{�{4�@ ���������������������������3���1163�>6 ��;;;?����?����@F  Nw�������������������������������3 fó���{�����{�?;B�``�c��������������������������s�??��1cc;@F�a���?�������?��>  �s��������������������������n6�?�3<43`6K9{��?����;��3�@ Bs�{����������������������������Nddd;C334�@Nc�������;{�� +C3s��������������������������d `B a6� 4�;;���{?{K��;a  g�3�{�������������������������   @ �C33�34 �a㷻�������;;4k� C?�s7��������������������������N@ `C�33�6 F�i;����{{;;����p ?�������������������������������FD@   ;3�ac� c�������a9;C3� s33��?������������������������Ld   c333@�;?���{;;�;do3� g�33���������������������������@L@ @�3c;C�� c泳����fFG�? C;6;7��������������������������Ld` F 3i;330 �Ci;���d���?1?@�4DF����������������������������FL  �@;333� F�;?{�<6�Ff �3c�36Bc3?����������������������������@d 33;3334 kc��93�f�@B;�?6D�;7?3�����������������������I��N �;;13� d���6�nB@�sc;c?1��4g���������������������`A� 3313�3 6C�6���KF@ ?;44333;s�?�7����������������������i��4��;3;3@n>�����n `33k0�1437��47������������������������ 337�33`hd3Ck;���� @ �;la�sk;;13�6f43����������������������99q��3�7;`�;;>c @` ;14C;;73s3?�CfC������������������������7�3334  K6����@ �33``1��?3���4f6f?��������������������4N;033�3;;{4$#k;;;D k  14FC�?�397;��6FfFO���������������������1�937?773�B �;9f` �  ��F�@����37��sdCfo���������������������;03�;s���3,` C���  �0 ����@ ?{s�93��6d?�����������������������3s�777?F��n64   7O����@ ��3?�?�6`F�������������������������;3����4$f�l`d��������FO���37���3�o��������������������������s1{�������C��k��������������;��������������������������������?��������K������������������������������������������������������������������������������������������������������