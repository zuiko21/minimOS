�����������������9���������������������������w������������������������������y?��D����La�?1��������������w�w���������������������������������;����tDI����������������������������������������������������C�K�9�d�;�?�����������s?w��������������������������9?9{���1�y�D�a�C�������������77??�������������������������9��������ƹ3��dDN�1�}���������==7���������������������������?9�����K9?�DL9?�������������w�3�s�������������������������;��9��3�Ɠ��?�������������{�?�����������������������q�?���;��K�1�iA������������������91�s�����������������������9�9�499���1��FAa��=�������?13����������������������3����K���99K;F��DN��������������s7��������?���������������4�9<c���3�9dD�AK����������;9A1;���������������������?1��;��a��9���D d��;��������<;w{������s�?��������������9�Ա���4ē�3���<dDD?����������;9C�w�����7?�������������1�A�96�aa�����L$�Ia�_��������t1<7��������1������???�?��?ә1�A�9D��?{���DFFL7�������������[?�������1?��{���{S���1��D�K�L��{��NDC��?������s�3��������{s��11?��y�99a�Fa9<d9�{;�??�cDDc���������F�7������w17��93[���9{���dD�A�;4D���?��{;ld������������1a1�w������9?��[�911�����s��LC@k�KD4�����dL;??�����1I977������717�����3?��94�L4I;�lF��?����9I���������������������3?�;q99a1;�;DFIc��K�O;?=��{y3�D19?��������w4ia77?���w��9����I11�;4{;4DAF�?;CAdC����������������{9A���?���3�;�4�Ô41�3={��LlaF��IND���������09��������41sw����7�94�4a����1;14DF�31�aFK?������?�������q��Ó����������o��IaiD9CC;��DC�a��A��i�����{{�K?s����3CAa?W����s9C�9Ki;9<11�DFC>1G����������������w�<N?{����31�a���a�C�9a�䱳;��;i��{��7��A��������4�CA����7����1�C�1�6�����KA;����y?�?q9;�4�9w����wD4�s�������3�C��K9ai1C�a4CA`Ĵ3󳳱{�{����9;���;9K;{�����44�Da�����7���1��I4�CKC�F�D��=1;3{��1C�����1�����{�{4�9��{s1C?3111�93i4��14KDdFK���;�{��;�����DKs{��w71AFD�����i?99;3CC��AlL1��[�;9��?4N=��;Da������;S�D��NC{������4�1��9;3���Kla��s�91��?�C����@D;1?{s�a�CD4A�����4�?�[�s���;ӷ��`AF?31A1FA1�4Dd@G��������ACI4��;�������I?����}?{��;�[�ID᳓IF@DLC?��C@@L??�0D?��1�1�9F��Ia4A������d����������?��FD1�dC�9i`DL??�D������[�S�1�DA4�C�������vI?�_������?���D @�91�KFC���DC������4D;��9�y;A�i14������C����?���=?�����@ i393;>DD?��>C?�����@�y��y�dDFA����C������D?�����{�������  C;���4  @D;��3�{??��@g�9991��IC1{s�������C���������������  ��3@ @  ䷿���1������@�ӱ�A`Dl3�����{��D?��������������@ g?4 dd���������0C�m��D@d1������w��L?������������� I��I;��1������������=����4iK�����{A��?�4��������������DG;�d��3�39����?�������=<9��{���y�?�47��q��4��������������@���;{3����;�����{����=��{=�������y����O��7i�������������DDC�?�����;�����7?�?������������������3��C��3�4C���������������A7�?{93C���{���������������������?��?��1{����������������B������9�_?�����=??��������;_�������9�����K�4D���������������F��??�{�3����D�??��������������������{C��A1d��������������� C;{���{�����{���C�?���������9�����������D��D�4L��������������DL{q?;{�i9?�?��D�{���������������������yd�d������{��������a7�;�{��1C������d����������������������C��dD����������������Lk��7�{sO�y{��{A�?����?���������������I��CLD����������������?�;�4;??7�{�FA3�����������������y��A�3LFD�����������������K;3�5���;4���d��{�����������������?��=<DD����������������4�����4�4���6�a����������������������A1FD����������������A;;��1C9FDii?�{1D���������������������{��KD�N@����������������;���;3I3��D3;��d;���=����������?������4�@D������������������;S�91d��6D��3������������������������1d�D��������������������94<fA;1��;;{�1;��������������{�����93��B��������������������;CD1�3�14��߷��������������������@DD�����}����������������dFA�1K?�����[��?����?����������Ddl������������������{DFLd<dDN;��;;??�{�����������������5;��������������������9idDDFDDN3���C[�?�=����9���������=�������?��������������������3d�k;;3?{���?����󛱱���������{[[������������������������a�D;4�?��39s�3����9��������󽿿�������������������9���=�1�694���i<��?���1�?�������������׽�?�������������������������4>C;���{7i���IK�;�������y��{�[�[��������������1��?��{�<443ii�����K4���{AL����������yy�����[�����߿������?����3K3������{�94O����������?��������������������������9������;�cCC�3���;��C0���3��������������񵿿�?��������[������������<<91�[3�9;I�;���?����3�������{��������_������{�����?�����CCK1��{{9��K�3�<�����?����������[9�׿����߷������;���������;31��y1@�;?9�������y?�������14�������������?�=�{;?���16C�93�33�F����3�󷗿���{�������䖔������[�������{����I�0D����1CI@���3������3�����������i1941�������������=���?1K�NCa���cad��1�=�������������������KL�����?�����?���������4�Al4������;󿳿7�������������1�iA4������?�����������=����dca�d<1cD I?�4�����}?��������������1a4������������{����������{���C��F��C�a�����?������������������d�����;991���3=�9;���ۛdcicDF@F���D;�������������������1idA�;993�1�����D��������99<IFKD<dDDA��L�?1����������������1K��;1�i�;[�?;�����4D1D<DDddFD��C�4K�������������������C1���>9kKC�?���������ۖDD��FFFL@KK�����{��11��������������9���6�a�1�9}=�?��?�����AA��FD�������;�O��?��������������������43�3����K������NiddND�0A4FA�����������������������3�13i11k6�9����?�?������ DAdDdC7@ �K�[�;��O����������������������;k13�?;�{�?������� F�FD��  KCӿ۟���?������?���������13�331�Cc��{�;�?����� F�D���@ �F��O���?����������������Dd11���1��13���;ӿ������9@F�C�4  ��A?������������3������{��LK��361�96[��@9�{�1���� DF� 	�;�����������1?�����������<CD1c�93�a31��������� ?��DDa�D�@C4M1��[3��?��1��3���������D<d313�43��3?��;�1 ����C@ND��1�D K99����������������������L31�aai<1A�����@ i�����D� 1K�����ӿ������=����������d1��C�C45�=3���  ����4 D���d@�����������������������FDD��13KCCC�c�󓿓@D��������D@[���K�������������������D�1��3i3IcCC�1�����9��4@F��F k��������[�����������������@@D;61143KCK6��L=3K��A����3 �dC��q�9�I�9������������������� a�ic�4444A�a�����{�i�{�@A�;@	��D �?���ۓ������������������4Ca3Ĵ446aa7��3���C��4F A9`�4co���?�1�����������?��������3<3�AcC��A���ѷC��99���d@ �a@N�q������?��������������3<16�1d�CA;��9;�߳���@� 	��NF@DDC���?����������������11C��CF�D<Fq9�������d@@{�D�6K�����O���{�����������������<<D�IdiDd�ۛ���;��D` �D��FN��C[1��Oy�����9�������������1C�D4iFD��@O��=��qI���DD FK?�1Lc���D�D�����?��3�������������kID4i�����0 K�|C������DDI���DDI���O����;�9��3A���������������DO������ �i�����4a�仿����O���������������������������a�� ������ �[������I1���K��;����a������������������� ?���O�@ 	�������{{@@�K����ID������=񱱐?������������������4 ��߱@y  ӵ�?��1�D�[�?<4L�����D;��������������������4�����4 C@  ��������dL{�A�����?������������������������@	���D@     ;������1���9������K�����D���������3�������������t O��D`     I1�����4K����ӗ�4����t K�tK�4����w��?�������?�� ���4L      C�����;?�I����9;�����0DA��9�9����{������������� ߱1�d@     �1�������41A1q�AA����@D�1���C���7�������������@K�4�D�    ?���ӿ�[@O� KD9D@�����K�C��1������������������K�D�I?�   �1�߿����@�0 �� ����t��DD�������s���������������A4FK��   ���?q=���4?��O��a9�����C�K�;����������s�������{���A@ D9��   ��?�6��6O�D@������6D@D��1���?���������������F D  I��   �ۙ�D���O4K��?9������Di��I{{=;����������������