���������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}��� ����UUUUUUUUZ���������"""""""""������������������wwwwwwwww}   ����� UUUUUP  
�
������   """"""������������������wwwwwwww    ��   UU  P    

��       """"""������������������wwwwwwwww}� ���� �P U       ��       """""""������������������wwwwwwwww}�  ��� �UP U    
� ��       """""""������������������wwwwwwwww}�� �  �UP     
���� �    """""""������������������wwwwwwww  ��  �  �UP      ��
� �   """""""������������������wwwwww   ��  �   �U   P    
���
�   """"""""������������������wwwwwww  }��  �        UP     ��
�   """"""""������������������wwwwwwp  }��  �        UUU    
�
�  """"""""������������������wwwwww   �   �        UUUU    �
�  �""""""""������������������wwwwww       �       UUU    �
�  �"""""""""������������������wwwwww       �       PUP    ���� �"""""""""������������������wwwwwwp      ���      UP       ���� �"""""""""������������������wwwwwww     ���     UUPU     
���� �"""""""""������������������wwwwwwww   �����   UUUPUU   
���     """"""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""�      ������ ���   www  w}����  ���UUU   UUZ��  
�  """"     ���   � ��   �        p    ���    UUU         
��   ""      ���   �����  ��   wp  www      ��      UUP  UZ�    ��  ""       ��  �����  �  �wp  www     �     UP  UZ�    ��  "    "" ��  �����  � �wp  www     �     UP  UZ�    
�  "    """ ��  �����    ��wp  www  �   �  �   UP  UZ�  � 
�  "   """��  �����     �wp  ww  }�   �  ��   UP  Z�  
  �  "   "   ���  �����     �wp  ww  }�   �  ��   UP  Z�  
  �  "   "    ��  ������      �wp  wwp }    �� �    UP  Z�  
� 
 "   "   ��  ������  �  wp  wwp p    �� �    UP  Z�   � 
 "    "  ��  ������   �  wp  wwp     ��     UP  Z�   ��  "    "  ��   �����   ��  wp   wwp     ��     UP   Z�   ��  ""       ���������   ��  p   wwp    ���    UUP   Z�   ��  ""       ��  �����   ��      wp    ����    UUU    
�   
�� """     ��    ����    �           ����   �UUUU         
��  """   "���  �������� ���  wwwwwww}���������UUU  UUUZ���� 
���"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������wwwwwwwww}���������UUUUUUUUZ���������"""""""""������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ������������������         
���������        ���������         ��������������������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@�����������                              @H@H@H@H@H@O�����������(�(�(�(�(�(�@ @ @ @ @ @   @ @@@@@ @ @ @ @�����������                            �@�@�@�@�@�O����������� ( ( ( ( ( �@�@�@�@�@�@@ @@�@�@�@�@�@�@�@