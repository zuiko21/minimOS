@@@@@@@@@@@@@@D@@@DDDDDD@   DDDDDDDDNDDNDDDDDDDDDDDDDDDDDDD@@D ������@@@@@���lF����D��D��������NNNNNNNNNNN@�@�@@H@��J@�,J@�@DF@@D@     @D@�LDDD�DLlNDNNDNND�ND�DDDDDDDHD $�$@@@D@d��LN@ @@@@@l lDdhlld��Dd��D��DND�ND������� D@@@@H@�$�@@@@@@@d�     @LDDDNDD��DLlDD��ND�NDDDDDDD@N @@`�D@D���lDD @NLDDd���D��LlldF��LFD�ND������� D�@�@D$�@D `@B@D���       `@�DDNNDLd�D��dLF��ND�DFLDDDD@� D @@`�`@��@D$@�DD@ @@@@ DNNNDDNF�lllF��dND�ND���d��� @`D L, D@�H@�d�� @   �D@d@DNNDLF�DDlFD��ND�NDLd�DDD@` `@@@@@D�@D$@D@�FL   @@L @ NNDD�dLd��F��lF��ND�d�Llll@ �D$�D$HD��LD @�DN@d @�DNNLLd�DF�dLF�dNDlD�Ld�DD@ �D@�@�J@@�@@L @@h@`D�`    Dl���@�`��DFFDlllF���NLd��ld�Ld��@ `@�D@�d  @lÙ;Ll@HD�DD�����D�lFDLdF�dF�Ld�DD  D@D�@@�@`�`@@@ �  F������d�dDNDdDldlF��d��lNLddDd��@@�@� @B�@,D�Dd�B@F@@ D�K����D�NDlLlDLF�lD�Ld�Dd����DDd  @@@@B@D D Ā �L @@@BF�;;���dld�F�FD��lF�ld�Ld��ddDB��� @D$� H@�B@`   DL;��y;��DH@D�F��DF�lF�Ld�Ldd����DDFD$�@@D��$@$�   @ d�ó���{9JF�d�dLlLlF�ldDDDLDddDNNNL@ �@�@@@@B$ @�@@�@ @ D�N99������L@D�LLd�dF�lDLNNNFNLNNDD�d @@@D��$�@H@�@D� D @@ @�diK�9�����dND�FLF��DDL$dDD���d�NNF� @@`@@@@@   L �Ʊ������4�NDND��DFF��LLllddd�D�DlF @�����B@`�@@�  @ @ D�㛳�����D�D�dllL@DLLd�D�LNNNNNND�@ F@F@@@@@`@�H @ @  �In�������F�LLD�$lldd�F�D�D�dDDD�D @H HHD$@@@  @FNI;�;��;�@NLD�FNF��FLLllLllNNNNNNLl d@$�H@  @  d�����9FND��lFNLF�DFFDFDDD�d�FD @�@B$�L�  @ BDƛI9����9�@NLD�dlF�D��LllLlLllllNF��@ D@@@F@@@B@@ @@L @   @FL<<����;�;�F�LLDlF�DF�D��F�D�DFD�lD @B�D$ HH@�@HD, @  @@��KK9�;��9�`�D��F�llLlLNFLlLLlllNF�N � B@HD@@@@@@B�@B@@    �BLi��9�{ۻ;@ND�dD���D�FFD��DddDD�DlD� @@@�@ @@�@@D   @ @BDFKI������D�LLldKNFNLllFLlLNNNLlF�F@ �@H@@�,@D   @  ��Dk���;;�Ld�D��d��d�F��F�D�DdF�D�@ D@@ @H@�@�`HD @ @@ @F�@D�;9;��@dLD�dNNFNLllFLlLNLNNLlld @�H @D� L @  @@L;�d���;@@LdlD��D��FDD��DddFD�FDF�@ d @@H@� @B@�@L    @  @d��DóidÛ@d��FDNNFNLllFLlLNLlllNDl@@�  @ @@@ ��I��N>D �dlLNId��d�F��F�D�DDF�lD@ F @@@ �`H$    � NDK;DỼ@@d��ddF�NFLllND�LNLlllF�� @�@@�  D  @@BH@@  D�@�dN@ �dd���LDLFDFDND�dFD�DlFD@ D L� @@@@H@JD   @D��Fƻ@K��DL;��FLNF��������LNLlllF��
@@D @  @   @ A��i�A�dN�K@ �dlLFA�LdNDLDdNFD�DDF�dD@ @�  @ @HJ@h@D @ @@ NK�Ļ�N��� @D��dlNF��������LNLlllNLN@@L @@@�@� @  @@l9<;9d�9���@�d���lLDdDdDdFD�dFDDDdFD   D �$ L@`@H@ @@  NK�ɴ�L;�9k� LDFFLFF��������LLLlllLLlDDh@@@@@D @@� @   A䛳�lD��K��@dllLFLlDLDLFLdld�d�D�d�D  �� H,@@H@@  @li;��F�9�;����dd����������LFLNNFLD��@F@@@@@D`@@� @   @@D��4NN��;�1 FFFF��lFDFDFDdFF�LFDDlFND  @ @HD@h@H` @@ �K9�DD��;�����NLF���������Ld�����D�@�@`BHD� �@D @   D䱻��K�;��@DddNDFLdLlDlFLdldNFLFDF�D@  `@@ @@D@H@�  @KK��d�C������D����F��d�D�D�D�lLlLN @D�D�@@D @@$D    @L99d�K�9���FDLlDdLD�DNLd�F�D�d�dDdd @@ �H@D��@  @@   d�@�I;��;@F���F��F�NNDd�LLLLLFLNLLL @B�@ND@@@D BDH @   LN LF�<;��DdDF�FD�lDD��NFFFFFLF�d�d D@ ,� `@��  @  @Hd� ��99� LLllDlND���LdD������lFLD�  $@@@@@�@`@D@@      NLD @LN�@�dD�NDd�FDLFLlDldldd�lFNF@ `@�@@@@�@@@�$� @@@   D�@ K�I9���LD��LLld��F�D�D��LF�D� @@�d�@@     D�LLDL��F���DLF�FD��D�dF�F�F�FLF�d�d  @ �@@`�@$� @  @ @FK;�LNLdlDLNdLNNLlDlLLD��lDLDL`DD$�@J@  H@  @@�@LLN�F��DNFLDldlNFDDF�lDddldd�ld�� H@`@H@@@D ��  @ �� ñ��Ļ�D�F�D�F�����lF����LFLD�FDH@�Ƅ @  @@@L   K@@D����@F�F�D�F�FNDKlF�FFFF�LF�F��  ` @B@@�� @ @@ K<DlDlD�9<lDLld���K�DlDlLlLDNlDLFD @D@$@`@ @@@  HiFHD�˱˴DldlN���F��NDlDd�dh�ldlND @l  @ @� @�  @@ N�dF�9;1�L@�D�K9��L�D����LLDK�D��D � @@D�  @�L @ FF���N���@ddNNLi�?�d�FDFLdd�D�FD� @N@@ @@ `� @F@ NDLll19kDĄ��û����ND����LLDK�LLND @@@�@@@@ ��@@ @  @@@D�d����� FDD�l9���?D�NDlDd�FNFFF�N  @ �@H@   @@@�@ HK�9�9<dD���LN�����ND�F��LL@N���lD@ @ @@H�@`@ @FF�9����dDDd�k���D�F�FLdd�A�dlD� @`D @  @`�`@ D ��D @li��9dLLlL<��9���NLlD��LLDl���ND ���h@  @@�@@@�@� i @@D���@@FBD�ṳ��DFD�Dd�d`ıFD�N @@ d @  @ H @@@HF@l@�L�������iik���<llFNLDLL�D�Lldd @ l@D@@ @ @@��d$@�FNO� `@lCN�����D�LD�NFFBF��D�� @@D �   � Hd@�@��� @D���D@l����;y�ND�ld�����d�ld  � �   @ @ N �DHD�dN�@�@@D�K��;��;DlD�LddL`D��lFL @`@d @ � @ L$B@@A O�`$K��F��KN������LF�Ld��FD�lF��  L @�  @ @� D����@DHF���� @@D�i�;����Ld�FD��L;��dD@@ FD$@ @   @H@@�@@@��>,K�L�`D @F����9����D��lLNFD�4NLN  @� �@ @ @@@@ @@d`d���Dl��C�Fl<9���������DF�d�L@K�LdF� d HD     `D � DD F�Ļ@Ɠ����;y���lllD�NF������d@ D  @@ @FD��NĴ�C���ii˱������LD�F�ND�@NF�Ld� @ F D@  @    �@@@�,@�l�D�9``@�ƛ;������dlllD�ND�����NF @��� @@@B @Dkd�lKKNC˴L9;������D���DDld�NDD��F�L @�@       @@B@ @@HD�K@�LF����a�BF˖���۳�NDllllF�ND��NLdld@ F@`@@ �@�D�@�NF�ilnN��DN9������INDD�F�ND�DNDdLD� � L  @     @@@F @@@DľDLF�F�i<� D䶛�۽9��dllllD�Ld��N��NF  FD @@@@@@ L D� �FLl�N��DK;����Dd��DFD�D�Ld�FLdL @@� �  @      D �@ @D@dKDLdFNC����Dồ���lNNLll�NNF��DNLd�� D @ @@L@ LHKNF��NN��Kỳ������Dd�DNDD�FLNĶLlD  ` @ @  @ @ `@B@,F	�D�d�9l�D�����9DFNNLd��NN@lN9;��Dl F�@   @ @@�D�@�@@@F��d��a�1��I9;���N��LF�LD�Dƻ���LiF @ @�@@@ @ �@ @@`@@d ��D���dlƖ��DK;����LDlld�ld�NNDi99�F�� @H@@   @  D @,�@D�lF��ii1d���?�?9d��F�LF�ND� D�����Ld@ `@ @@ @@@@�` BD��lF��NLK������LDllF�Ld�NNNNDld�F�L @H@ @     @ @@@@D L@IlD�Ll�i鳓���D�NF�lD�LD�D��떜FLd�   @@ @@@@@ @�@�@$N�N4�llLF��;���LD�lF�NF�LdFNC�f��ND@@@@Ā@     @@� @@@�@�H�D�KF��d�K9;���Ld�lF�ND�Ld���I;��ND�  ` @@@@@@ BD @@h@D�ld�l@Ld;K�����ND�ld�ND�LlFD�FD�ND       � D @ @@D @DNLNK@D��;���4F�NND�D�ND�DlƓ���LdN  D@@   H �@@�,�,��kD�@@�����?��NDd�llND�LlFLi9lNF�D @@ �     @@@@`@@@DKC����KK=�dNDlNLD�D�LdFLd���d�d�  @   @@@@@@@� �lKld B�乻��D�F�LdldLd����La�NLlND @@@@     �@H@@FD �@KƖ��D@�K;K�D�F�LF��LdFLlF��D�F�N@  @L   $  ��liN @FK����4�ldLd�dND���F���lIld @@`      @@�@@@@@F���@���LDNF�lND�LdNLdLa�d�D�  @�@  @B@@��  @�KN@@DC����FF�LF��ld�LD� DD�LdLd @@` @@     @�@�@@@�@L`D䴴 @�99�LLF@DDF�Ld�NDD��llNFL@ @@  @@@@@� @@` @�FKKD H@�@F@;���FFĆ���FD�LD��a�FD�d  @ @@     @ @D, @@@@H@  ����D �������DdFF��NF�DND�i�NF�  �  D �@ `�,$FKK@H@D` DL;�DDddNLLLDdDDD��@aKA�lF@@@ @     @@@@@D�@@DH l<`@`�$ K�NNL@�FFNLllldD�Γ�LDl   @@@@@ @@ @D NK@�D�@@�D�DDF�@���D�D�D��FCľF�D@@  @@     H@ @@FH D`�F @@C�� B @��F���D�ddd�F�F�DF�L;�l�  @@  @@H �`@  NK@F�F�DFLDDDlDLLLDLLLLLlD��F�D    @ @ H @@@@@@�D @@i9 @$ �HFNNNDl`ddlddddd�`K��D� @ @@ @@ � @ @�@d�@ N� H@L@@@DdDDD�����������LND�>ND@ @  @  @@ @@ @L�@� D @D�@ � BL��F���FDFFFFFLFFLFD�䳛D� @ @@  � @@@$�`  K@ @@D@@D�DlDDD��������lLd�ĻIi;ND @  @  @  H@ �@�@@@�$�@@`�dDlllddFFNFFF�d�Dd���KDN @ @@ @@ @� @ L �D,d@�DDD����D���lFNLD�i<�D@ @     @@$�d�@d  @HH@@@BD$���dddllddlFLDFN;��� @ @@ @�@H@ @@@@�@@ H@ LD`DD�LLDD�����D������ĳ�<D @@     @@ @@�D @J D$D�dlldlddd�NFDdDDd�;���N @ @@ @@@ @ @�$ H�@@HD @NDHL@@NLDD�D���LD������N����D@@H    @ @@@@@J@�  H@HBDND���F�FND��DldLF@9���� @@@� @@ @@� B@@H@@@@B@H@��`D��NDDLLD��NDF����d�F�9�ND@@  @��@  D @@@�@@d @@F@@DdDDNNFF�Ld�NLDdlD�d˱���N @@@ @ @ H@@@@@@@H �BL �ND��L,nDD��Ld�ND���F�LNA��i<D@ @�  @@ ��@@@$ @@D,@DB@LDKN�lld�D�lFD��LFDlla��� � @�@@  @ � @@@@�$@ �� @lNN�DFF�LlNF�lNND�d��F�ÖD