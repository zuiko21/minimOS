                                                                                                                                                                                                                                                     """              UU           �������           wwwwp        �������        """             UUUU          �������           wwwwp        �������        """"             UUUUUP         �������           wwwwwp        �������       """"            UUUUUU         �������           ww wp        ���            "" ""            UUUUUUUP           ���          wp wp        ��            "" ""            UUP UUUP           ���           wp wp        �����         "  ""            UU  UUP          ���           ww  wp        ������         "  ""            P   UUU          ����           ww  wp       �������           ""                 UU         �����         wp  wp       ��  ����          ""                 UU         ������         wp  wp       ��   ���          ""                 UU            ���         ww   wp             ��          ""                 UUU            ���        ww   wp              ��          ""                UUP             ���       ww   wp              ���         ""                UUUP             ���       wwwwwwwwp             ��         ""               UUUP             ��       wwwwwwwwp             ��         ""               UUUU              ��        wwwwwwwwp             ��        ""              UUUP              ���             wp              ���        ""              UUUU               ���             wp              ��         """"            UUUP              ���             wp             ��        """"            UUUU               ����             wp        �    ���       """"""          UUUP              ����              wp        ��  ����     """"""""""        UUUUUUUU        �������              wp       �������      """"""""""        UUUUUUUU        �������              wp       �������      """"""""""        UUUUUUUU        ������               wp        ������       """"""""""        UUUUUUUU        �����                wp         ����                                                                                                                                                                                                                                                                                                                                       ���������������������������������������������������������������������������������������������������������������������������������������������������������������������  ���������������  �����������       ������������     ��������       ��������    ��������������    ����������       �����������     �������        ��������    �������������     ���������       �����������     �������        �������     �������������      ���������       ����������      �������        �������     ������������       ��������       ����������      �������       ������      ������������        ��������       �����������  �  �������     ���������      ������������        �����������   �����������  �  �������      ��������     ������������  �    ����������    �����������   ��  �������       �������  �   ������������  ���   ���������    ����������   ��  ������        ��������   ����������������   ��������      ����������  ��  ������         ���������   �����������������   ��������      ���������  ��  ������   ��    ���������   �����������������   �������       ��������   ���  ������  ���   ��������   �����������������   �����������    ��������   ���  �������������  ��������   ����������������    �������������   �������         �������������   ��������   ����������������    �������������   �������         ������������   ��������   ���������������     �������������   �������         ������������   ��������   ���������������    �������������   �������         ������������   ��������   �������������     ��������������   �������         �������������   ��������   �������������    ��������������   �������������  �������������  �������     ������������     ��������������    ��������������  ������� ����   ������       �����������    �������������     ��������������  �������  ��    �����           ��������        ��������       ��������������  �������        �����           �������        �������       ��������������  ������        �����           �������        �������       ���������������  ������        ������           �������        �������      ���������������  �������      ������           �������        �������     ����������������  �������      �������           ��������        ��������    �����������������  ���������    ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������