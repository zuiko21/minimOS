                     DDDDD     DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD                     DDDDD     DDDDDDDDDDDDDDDDDDDDDDDDDDDDDDD                     DDDD@     D@DDDDDDDDDDDDDDDDDDDDDDDDDDDDD                     DDD@         DDDDDDDDDDDDDDDDDDDDDDDDDDDDD                     DDD@       @ DDDDDDDDDDDDDDDDDDDDDDDDDDDD                     DDD       @  DDDDDDDDDDDDDDDDDDDDDDDDDDDDD                     DDD       @  DDDDDDDDDDDDDDDDDDDDDDDDDDDD                     DDD           DDDDDDDDDDDDDDDDDDDDDDDDDDDD                     DDD           DDDDDDDDDDDDDDDDDDDDDDDDDDDD                     DD@     D     DDDDDDDDDDDDDDDDDDDDDDDDDD     @               DD@     DDD@    DDDDDDDDDDDDDDDDDDDDDDDDDD                     DD     DADD  @DDDDDDDDDDDDDDDDDDDDDDDDDD     @               D@     ADDD DDDDDDDDDDDDDDDDDDDDDDDDDD                     D     ADD@DDDDDDDDDDDDDDDDDDDDDDDDD                     D     DADD@DDDDDDDDDDDDDDDDDDDDDDDDD                     @      DA�D@DDDDDDDDDDDDDDDDDDDDDDDDD                     @     DA�D@DDDDDDDDDDDDDDDDDDDDDDDDD                        @  DA�D@DDDDDDDDDDDDDDDDDDDDDDDDD                        @  DDA��D@DDDDDDDDDDDDDDDDDDDDDDDDD                        @  DD���D@DDDDDDDDDDDDDDDDDDDDDDDDD                           DDA� DDDDDDDDDDDDDDDDDDDDDDDDDD                          DA� DDDDDDDDDDDDDDDDDDDDDDDDD                           DA DDDDDDDDDDDDDDDDDDDDDDDDD                           DA DDDDDDDDDDDDDDDDDDDDDDDDDD         @                 DA DDDDDDDDDDDDDDDDDDDDDDDDDD         @                 D DDDDDDDDDDDDDDDDDDDDDDDDDD                           DA DDDDDDDDDDDDDDDDDDDDDDDDDD                          D DDDDDDDDDDDDDDDDDDDDDDDDD                           DDA DDDDDDDDDDDDDDDDDDDDDDDDD                         @D DDDDDDDDDDDDDDDDDDDDDDDDD                          A  DDDDDDDDDDDDDDDDDDDDDDDDD                          D@DA DDDDDDDDDDDDDDDDDDDDDDDDD                            DDDD DDDDDDDDDDDDDDDDDDDDDDDDD                        D   DD@A  DDDDDDDDDDDDDDDDDDDDDDDDD                        @ @A@DD  DDDDDDDDDDDDDDDDDDDDDDDDD                         D@D  DDDDDDDDDDDDDDDDDDDDDDDDD                        AAD@  DDDDDDDDDDDDDDDDDDDDDDDDD                        ADDA DDDDDDDDDDDDDDDDDDDDDDDDD                        AD DDDDDDDDDDDDDDDDDDDDDDDDD                         DDD DDDDDDDDDDDDDDDDDDDDDDDDD                         DDD DDDDDDDDDDDDDDDDDDDDDDDDD                        DDD DDDDDDDDDDDDDDDDDDDDDDDDD                         DDD DDDDDDDDDDDDDDDDDDDDDDDDDD                          D D DDDDDDDDDDDDDDDDDDDDDDDDDD      @                   DD DDDDDDDDDDDDDDDDDDDDDDDDDD      @            @      AA DDDDDDDDDDDDDDDDDDDDDDDDD    @ @                   A@DA DDDDDDDDDDDDDDDDDDDDDDDDD    @ @                   DA@ DDDDDDDDDDDDDDDDDDDDDDDDD    @ @                    DD   DDDDDDDDDDDDDDDDDDDDDDDDDD    @ @                    DD   D DDDDDDDDDDDDDDDDDDDDDDDDDD    @ @                   @D@  AA DDDDDDDDDDDDDDDDDDDDDDDDDD    @ @                   AD A@DDDDDDDDDDDDDDDDDDDDDDDDDD    @ @                   A DDA@DDDDDDDDDDDDDDDDDDDDDDDDDDD    @ @            @      A DD DDDDDDDDDDDDDDDDDDDDDDDDDDD    @ @            @      A@ DADDDDDDDDDDADDDDDDDDDDDDDDD    @ @                  @  DDDDDDDDDDDDDDDDDDDDDDDDDDDD    @ @                  DDDDDDDDDDA�DDDDDDDDDDDDDDD    @ @            @     D ADDA�DDDDDDDDDDDDDDD    @ @             @     DDDDD@DDAD�DDDDDDDDDDDDDDD    @               D      DDDDA DDDD�DDDDDDDDDDDDDDD      @             @      DDD DDDDADDDDDDDD@DDDDDDDD      D              @      D@ DDD�DDDDDDDD ADDDDDDD      D                   DD@ DDD�DDDDDDDDDDDDDDD    @ D              @@   DD  DDD�DDDDDDDDDDDDDDD    @ D               D @   D  DDDA�DDDDDDDDIDDDDDDD    @ D                A@   DA�   D@DA�DDDDDDDD@ADDDDDDD    @ D               @D   DO�   D AA��DDDDDDDDDADDDDDDD    @                 �    DD�   A��DDDDDDDDDDDDDDD    D                 D�@    D�D   �DDDDDDDDDDDDDDD    D                     A�@    D��DDDDDDDDDDDDDD    D D                 O�@  AD    A��DDDDDDD�DDDDDD     D                @� A   A��DDDDDDDDDDDDD                      @DD AD   A��DDDDDDDDDDDDD                      @D@DD   A��DDDDDDDDDDDDDDD                    @ D@DDA@  D���DDDDDDDDDAADDDDDD                    D DDDAA  D���DDDDDDDDDADDDDDDD                      DDAADA  D���DDDDDDDDDDDDDDDDDD                     @ ADDDDDA A����DDDDDDDDDDDDDDDDDD                     D ADDDDDDA A����DDDDDDDDDDDDDDDDDDD                     @DDDDD D��DDDDDDDDDDDDDDDDDDD                      @@DDDD@D��DDDDDDDDDDDDDDDDDDDD                   @   @ @DDAD��DDDDDDDDDDDDDDDDDDD                     D AD  DDA��DDDDDDDDDDA�DDDDDD                    @   ADDDDDDA��DDDDDDDDD@A�DDDDDD                      @ADDDDDADA��DDDDDDDDD@ADDDDDD                       @DDDDAD���DDDDDDDDDDDDDDDDDDDDD                     @  @DDDDDAA���DDDDDDDDDDDDDDDDDDDDDD                       @DDDDDD�DDDDDDDDDDDDDDDDDDDDD                          DDDDAD�DDDDDDDDDDDDDDDDDDDDDD    @                    DDDDDD@D��DDDDDDDDDDDDDADDDDDDDD    @                     DDDDD@ D�DDDDDDDDDDDDDADDDDDDDD     @                     DDDDD  ��DDDDDDDDDDDDDDDDDDDDD    @                     DDDDD   A�DDDDDDDDDDDDDDADDDDDDD     @                     DDDD   DADDDDDDDDDDDDDDDDDDDDDD     @                     DDD    DDDDDDDDDDDDDA�DDDDDDDD     @                     DDD@    ADDDDDDDDDDDDDD�DDDDDDDD     @                     DDA@   DDDDDDDDDDDDDDDDDDDDDD     @                    DD@     A@DDDDDDDDDDD@ DDDDDDDD     @                     DD      DDD@DDDDDDD@@DADDDDDDD                            DD     @DDDDDDDDDDDDD@DDDDDDD                            DA      DDDDDDDDDDDDDDDDDDDD                            DA        DDD DDDDDDDDDDDDDDDDD                            DA       ADDDDDDDDDDDDDDDDDDDDD                            D      DDDDDDDDDDDDDDDDDDDDD                                  @DDDDDDDDDDDDDDDADDDDD                            @       @DDDDDDDDDDDDDDDDDDDD                                    DDDDDDDDDDDDDDDDDADDDDD                                   @DDDDDDDDDDDDDDDADDDDDD                                   @DDDDDDDDDDDDDDDDADDDD                            @       @ DDDDDDDDDDDDDDDDAADDDD                                     DDDDDDDDDDDDDDDDADDDD                                      DDDDDDDDDDDDDDDDADDDDD                                  @  @DDDDDDDDDDDDDDDDAADDDD                                 D  DDDDDDDDDDDDDDDDDDDDD                                 D  @DDDDDDDDDDDDDDD A�DDDD                         @       @D  DDDDDDDDDDDDDDDDD ADDDD                                 @D  DDDDDDDDDDDDDDDDDD�DDDD                                  D   DDDDDDDDDDDDDDDDDDDDD                              @   @ @DDDDDDDDDDDDDDDDDDADDDDD                                 D@ DDDDDDDDDDDDDDDDDDDDADDDD