DDD�DDDDDDDDDLDDDD�NLd�@@@@D��LdNNKNKKKKKKKKKKKKKKNNNNNKKJNJFB����JN��F�����id��I���i<d�D�L4Ɣ�䴴������������4�1�lDDDD��LDDLd�D$�l@D,NLN �@HDINDNN�4�N;�������Ö���i�Ik���뤆��d�l$���B��d�NJFD��l�DB `@N�D���F�L��KKKKN���Ɩ�i��<L4DDND�D�LDF@�dLF�`�DLFLNLD�$�D�LL<ili<<ᴴ�����ll<<ikCl<F��h�NBD`hLlD��HlLd���<4�@H@@��LFC�ĴƖ�NKKKKNKKKƔ�C�ļaDBDLhLD�FDD�@dHBD��N@  `@Ll@lLiN������ᴴ����iid�<kFBĄ���BJD��LlD���Lla��@H@ hHB�D,@l<d�N��KK���ƖƖ����K��Ni�DB�Ƅ�JBF�lD�@�F@�iF� LL��KKÖNNi9iiiii��l<���DJL��dd`DLDlN@�dLd�F� H`@�d@NL$LDĴl<ll9a���������l<i�Ld��J F�����hFD�LdND�d�d� @lc���dHd�F������KKN�Ɩ�d�IkHDLJFDFB@D�HHd�L�LNIf@��Li��>��DHlKNIli���������l9l���F�@F
FĄ����F�LD�D�@�� L B@d��߱�N�D�d��ÖiKKKK��<nLd�9ND��d$LdHL@�D�F@���N@�F@N{��9���K���iin�Ö����ilC�a�KN� ��d(LH@Hd`�$�d��@�B� @�@d��������NAl;I斖���<<<<<<f�a�C�<��<DBDHDNF�@�D�LLdlNDld�@�D���������NƖ�KN<1�����NF�a�a�<�HJFJDL�B��Ą`N�L@,N���?����D�<<<c�����NKD�c�C�i��<BD�D�$�`HLD�D�D��F�$ D @FC��������<lNKĴ�<��d�L��i���il� d���HLd`�d�ldN��d@�iɿ��������D���<il��NFF�A�N�<�4�Ö�NH@HLNFFB��LHD�D�LLd  d FKc[�����D�lC���<<�C���KK�KK����dJDFB�FJF�D�N H H@B�˛���������FĴ�KId�NIk4�Aia��i��nKNJH`�D�`FFD�DLL@F�@@@ �NC���������HIa�NIkNiL�;�i��<<<������D�LNF��N�Ć@�  �l��������FNNᴴ��䖳K��C���l>KKND$N�DdHD@@�D�HFD@@$ llû��������Hi<kLd��ᶔ�����i<����IiiiHB�@LJNdNF�B�HN@h@ @FK����?����ND�>KIkiiCKC��KKKd����Dll$D@�DDHDF�@ H����y�������lil9Iii䴱������������(@�����L,lBF�ƄNB@� Ll;�=������@�����KNIkK��ia䴱��N<>D d�L$@dd@@d�@LD�D� B��D���{������nL9Il��Ö���iil9iKIiN�LdL,LhHNLH`��l� `�@@J@NN������FIf���ᴴ��ô��<6���Ɩ�����@H`dhN@@D$�LDDF�H`� �I������HF���������ı��i����������HdD�D�Ƅ��FNB�Ƅld@@ �N�D���{�@LKKNi;N�<<<<<><>KK@HHl`F
D@F@F��DLD@@� @`@��K�J��1���NKCƖ�������l������䔴K�FHDJHLHDdƆ�@@�� B��A��K�9@<9lii�����Ö��K9l<>kK�@LBD�DBD dDD@D� @Ą�@@@��K�l���F���Ɩ��Ö������䖖�䔴K�LBFĤhL,LBHD$�Ƅ`�$ @K��4a��A�[KKl<i9<<<9i<<1�KKKKKii�@�@L@Dd@`D�hLdLD �� `��F����dNA�@��KIF�����KKNL<�����ƖKKD��NhHHHHHL@D`L`h@@`D��n�i��K���@���i��<4�����NNH$L@@D$NL`�F�� @@I����A�{K��D��La�9i���䖔�<ilKI4����@��$�l(D��LLLd`�F�D �@�9��?�������K��KKKKiid������KK N�DHd�`BD��hl@� �BF�[{��y��F	l4�il<ii����Ɩ�KL<IA����HFDd�dHdF��d�@l@@������i�����HNA�l䱶��i4�����KikK@lhLD�$��DLd�$�@@� �@hD���KN�����@KNKCIl9ii���䶖�KIl><F��JDD��dd,ld�dL��� lA���F��[����iid����KKKKKKIl4�������;K@Bhl@N���@H`��l@`  H;9��LC�����,NNIdf������IKiNiNKF����F���FFD$��D`@�HhLJ@LĻ��i����Di�K�i<<<<1���ƴ�i9<9i<@@�@�@d����D���LdD @  K����K���߹HN�KD4Ɩ���Ɩ������d��Ɩà�@��FFF��B�L$��@@HL@�9��K���~FA���<9iiiKI<<l>���iiiD@�L@F�`hHHLDl@�L` $  F�;@DK���{�LN��1Ö����������NN�Ɠ�� ƄF���`hdlD� N  N LL,a�L,�;?���i����N�<kKLikF�L<I<il4���H`�HDN�DD�D��F�@ @H J  Dƛ@Lk����D�KLi�Il9iC��<c�䴖���iilhJD��B�$�N H@� @@D$��ihJD�?��i�����Ɩ���i4ƜlKliK��B��d@DNLld$` `��@�K���DK��K۔F�lC���9l<<<4�NC������iiJFL`ld�����@ĄD 
D����컿N;D�k��K���Ĵ�䖖ƖKKd�ᱴ���DDF���@�B��d `�K�@L3���I�@<D<a��ı䴱�Na��Ö�Id��NN@FllD�����@D@Ĥ@@�@���ND���9;il�NFNKK�<l<ll��l<����@�� ND@@D���BD��NH `HK��FDC�ۻ�C�I4��鱴����iiC�<<;��KN@DdNDNLh`DD��DF@@Hd���i��NInLN���K�N�Ɯi��K�������� L��@@D$L
$���`@N��DK����ƴĶ��?������<<a�IlL�KIlIiHlF�l,NHLL D���B@� �hD3���K;�INN1����������Na;���ᶖ Hl�D@`@`dL@KDND F̓������@NiC�Ii�����a����l9lL�NNIi@DDNHLHHHlN@H` HL,F<;�����Hd�L<�������ilF���F�KF��Ö�$�@d@dd@@@D`D��`D�ND듓����d����������ii>��iiL��iilii@@�D$�HHl � Ć�Dd��IhL@��C�����NKD������������i<KNF�������@ldFd@D$�BDHH@@d��L�9��DFL<ND�������a�����ğ4��iliiHh`�LHN �@@��dl@�������K�9y�NHF�Lk��������K<N?�id����DDnF�D�D��DK �l$D�9���d�id��;�����KKKIliiKd�9K�����`@��N��@@@����D�,�O�@��N������D���;�����������KKKI;��i<<<4 �F�FNL`hD D@HN��L��lDl9��$D�	d��������A���Ɣ��ûᖖ�KKKLƀ�BL L@��D`NDB@�L�D,llD���L,D˹�������KKNNiii��� `BDDnL �� @�F���hL$K��D�Fƛ�dFLA�������������䴴L��KKCƖ�BL�� �@F� @F @�BD$�$LK@���JLK��Ą�$k�;�������NNC�󴴼<<1 @@dNF��B(HlBL�FĆ�O�<D�?���@d@ě;߿������ᴴ���i��KKCÖ�@J$� ND DBd,hd�FD��K�N�K�HdN;ۿ����������NKIK;����<ia ld��@ hL@�D�D,ldlNL0D���F�l���������KN����L��Kia�Þ��$���dH`@ ��H@d�FL9����ÿ��dÿ��������䴱kKKK�o䖖���@@�@l$L`@
H`BHFDd`lF�L�NKK��;��$LK���������KN<iKK�k9il FL,@ @����JH@@FNDƹFƓ�;9�Ĥ�������ñ�ᴱ䖖�la�������H`�
L@ND @@�@BDF�����$�L<i9����@Nۿ�����K��KN<<KKK�Ö���� @H@NNDN� @�@���dFD�O��ƴ;�?�LC��������l<9i����ᴓ�l<><<1D�@@�dL$@ �,@@@��LN�K�<iK�9��?dl���������<<<<<����KD�NHd  @@@@HD,L,`d�d�D��䖴C�����ý�����������KKIi������L @�DĆLH`��@`D��D�LlD�FDƔ�9��4�;�������������inD䱳�K�KKK @�BL @@� B@@���`Hd�N��Ll;�9{�K�����CKKKK��N����a����@�@@�D@ @���@l@hD�$Ld�O�d�ñ������������˱���l<������>�(,JD( `@�LB�lDhd�$LD�<�99�9��������<9l�����ilD�����iiiiiH@DD�D@H �HF��N@���K����i��Ώ����C�Ö�����N�Ó;?�; �@�Dl , B�H@�D@FJD�F��K��L������<<9iii<4��9l;��3�����@L D�@@D�Ą�`�DN��F��Þ�9F��������KK�������ü9�K��KNHND�@�@@�B@$`@�d�@@D,�ļ;��䑿�����l����iiid<iC�9������B@@B�`B��@�����$H@FJJND99iai���?���A�Kiil<<�NÓ�9i>KKKK@��@�L� B@,@DDD,H`Ƅ�DDH�����D���������Ö����C�ii����������@�H@, �@d@FNN��KK�<;DNI;�����KI9iiil<���ƛi��ikNKKK@ @d�`�@@L$�Ll,HD�D@�91��D���������˖���9����ᴴ���BD�@�BB`HD@FFF��@��K���@��d;ۿ��iC��Ɯi������K�ᴴ���$,d$@@ Ƅ��Ƅ�D�$LF�9��@dē�?����li<iic�CN9�ÛKKKA@� FL`��D ��L@DNDJN HBI����LL,o����KÓ����<��Ɠ��;�N�����@�D�� D�J@D�,h`NFLDLl�9d�@FDL������KN1�C��lD�<�NKKKAH@`�D�$� �@DD�@�D��� @γ��DDLD����NLd����>��NdN���iiii�B�@D�l @Ĥ �BĆ�@�D�@N���DKK�J@�D�i����>LdNKC�in���Ki4����1 @�@@ @ @BLDlNNF ���Dd@@NDD���D�I<��ƞID�i;�˱����L$�F@B@H@�HD�@LD,LL@��i;�������K���l���l<A��KLN��4��䖓$ ���$N@d$�B�D����� hK��FHDH`LND���LFLA�Ė�4��D�������@HDd@@H�H@���@�D@@@D@D仴HdldFD��<d�L���iNkNKL��iiKi<>�@HB�@@h@LDhD$�����A����FNLl��I�d��Ɣ�����a�����ii@�B@ d,,@���H@,hd�@λ��D�FLF�Id�l��inKkili�����Ɩ@@h@�@�@@$D@�@��lllBL@C��D��Ld�$�ll<iC��Ƒ�Ɠ�K����Ô�D�@�D���HD��@��dFĻ`$Dld�d�LF�����l�iNN<KK����<<kN @`@,�@ @�BH@D�NLNN���F���H`L`�lIl<�n��Ô��;������9N���@�`@J@���DL@B@�d`@���Ld�Ld�LKF�KD����LllkNKO���<iF�B@@� @�JD@��B@�B���`Ą��F�D�@�F��NF��l<��KKiF���Ĵ����FD��H�@l �� ��`d@�,d@$d@�D�FD�Ll��Nil9lilKKl�۱�L�<��`@�F@hB@�@�LLH`LLLdDL@FĄLlllFNF�d��Ɩ������<4������KI@@ĆD� J@@�`JFL```Hh``HLN@�DFD��Ld�NIn<>��n�{��iᴶN@$��,H@B�D�D�����d��HB@��F���D,dƑa���������9d�K���;F��� @�����BH@@�@F�DdN@d�FJ@@��FF�DND������<i<i<>NIn1���KKiD�$@`F�B�@L$HD,D�dD��D��lLDlNC�IlikND����D����,�@�J@@@�D@lD@Ldd,D�H@��`d�FL@d��4��Ki�㖔������������K<@DF @@@@�������@HLF�`DLLFHLd��NL˴�D���Ɩ����i9N9����l������JD��� ��D�Fd�LF@HJF�HDlNLld�4�1�<<l9iK>�Ɣ�;�;�Cù�F�BD@F@�@H`�HDFLD�
@dLd���lFFLF�D��Ó���k���KC�A仓�d���