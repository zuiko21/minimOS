?��?�1C3�1@�334{11;�CDCO3��414DDC1C33133333333D07@C@�����D��@99�3��O?�3�49��dO�1?��DdA�O[4Iy9;49?a?F@3���;DK?d4KC�i43C��=�C;�?{;�14dFC;433�FD131�33 07@����1D?0�IyF14DK{{1�;3�1�?1��4dC�����DF@G��4;6D?F{�{��D��ƴ0D�D�1���3��?3�C4KDi;D134FDFK314�sD`3A�����;D4�A40 � �4KK[119;1;;{s�1�4Dd��DDd4O9;3�4��D`F��K��4�At 4�O;C;1�91�?;3���;?7�dO�4��47�dD�A�3d�?D�`�0A �����K9?��A�4�O��[���7�?3�4D�;@K�d4cD�C@C@@F�����C�{10�1��3��?�;��{��;K[1o���K@DiCD�d{F4DD0I����A���1� ��;vo�1�[��9?w��3�����;DD<44��7DC4DdDD0DC�?�A��A��D� ;�K��S��1�S�?G�1??4ᴴa��D��?K0D�F�@D�����;D��d4;?a�1C?�3�1��1��?;�?�����4K1�4t�4D 4@dG1dDFD�����D4����K��q��s;w��;��93;;�9;4�K;�D@K�DD{���D�C�FtD�9D{1�{{1����?;�{�?��3��3���C45��1D0CD4DD�{���3D�A�4�D� D4@������7�������?�����A���DCKD�A@DF@�����A���4�d��O?�����ay{�?{���?;;?��K4{�DLCD4@ D����F�134��C��t1?�;����1�;�?7���;{������1a�1�9Da�DD@DDF@����D?���	3�44�?���7?C����9�?��{�?�;����;@D@4@ @D�����444 I�1D;����=?��1���??{��?3��{�4��DF @@D`D@����3;3��D4@�;�;C��7��;�{�;;?��D��K����;D@DAD  D�F@�;1����;{�󱱱1�O3�s�?��;{W����;43�FCTd91;CK��D9DDDD=��3�=�����{���?��;�}?��{?�{���?���sCK�DC�D9�GKC  @@D�;�{3;y�s�???���1�����;����?���{��;C`D1��4DaD@Dd@A�?�{�����y���{y;;?����7�?�=����{{3�KD���D�AA 3@K;��;1�1;���??9�{��a��1;�3�{_󳷳��1C@�DA4KKD1F�4DOD���??����������991�1�3?��?;9?�y�������F�D@DDaD1@�DcK?F��C��������������{󳟷�����ױ3�;�O����4;9d`D`DDA���AKFK4C��D��?�����{��?����������{;{�{?��?�K��DDDD�C4DC�A?�O��������������?{������?�������1d�{4��;ADDa�aFK�C�A;?0A��?;����������������;����?��K��;?�� dD�AF4DDO�DK;@DId���9?�����w�{���?�����;?��1��@O9��?�;dDdIC��D�DA�D@ D�G�����������?�����3?������9s���������D`�DAD@��dD�@ A9{��������7���������I������?��3���tC;;D@4DD�D4�F�@ DN����������?��{�?�����9s���4;?����������F@D�DD4�14A�D@0A9?�����������?���������4��DDI����D�{D@?�D�DDLD�D�@ K@C�1������������?������7����1�@@C����� ��<FA@@DDF@��DI�����������{������4�����K4dFD�����3D;;A@KD4�D�d�t D@C��?�����������t@��������94�KC��;��FO�lDC�333cD IdD4��K@K�?��������{��{���0�������i;KAA��O<D;4FDO{{��3@C�@C�D@�O��������7�����v��4A9����3FC�{?�0 C�4dFC3�1193DD@���D����{�����{�������4�F4�aK���A?�K����4Di3�Ad�14�CFdD@DC4O�9y��������������41�9K���3�t�Ad�1��4C�4d�;;33�D�Ck KD?{9�����������������ND�4������Ay��;����?<F@I3�a�4di@?�4�����������������dd?�������1�	4����6DD��d@31��44FAf@�dG@����?����������4D?4���?A�C��s���0K�D@��91��iF��@6�;D ���������������?�d�4K����C�C�0����{F��FD33�3��4;0�;4��������������������@?�A�����I?KCA�?������;D{1�49a49931N�@������{��������?��K?4��;A��C;�I0���{3;�DC�9;;�K����Dm������9O����������O3������K�dDO����9{4F�3�1�;11d130pKD������������������?�o������C�@ ��?6��D1;3�d󔱳��y�0D?����LD����������K3��������A�	4DDD���;91�>A�7��D4CK<� D�9K�KD�@����������0?��?������C��4����;��K� A�;1�KDi?�?O�@@����I9@ ?���;?;{�;��3�D���kyC�������3�9;�@1�aCFC��@@��D@DDDDDDDK��?��D@@D4;�p{1�����9d3�����KF�A��9?3��DA����DD   D@@���DDDDK��?����??{�A���;��14dFA1���{d K�<FK@DD @@D ���3@@C?��0���;?��4C?��I�����DC4t���D�C�dI�D D@@D@D �{�D@D d1�p�������1;�����9�FDC���q;�DD�LID<DD DD@��t4DD@a;������4��3���{��ɹ��>D44t����<F��FD@@@  @@?�?��D@Dd4��O���?�����񴑹��A3���1I@DDIADD@D@D@@��?�@DDCA�����9?����?�����������A�i?;NF DDL4��DD@@@@D@o��4�D@@Dd��9������������������ə��CD1�C91dDD�D@@D  D  O�;10D@DID������D�����������9�DLKC3�D1��DFI�NDD@@@@@ D D@O���@C 4���������������<9�D���K�49d DaDD�DDD@@ @ �;4ADDC���ɑ������� ��?���D���D�Dda4KDD@DF�DD@@@ @@@ @����D Dd@I��������O��� ���������<A�A�4D;;4DDDD�D@D@�;9I@ DDc���9�����D@�����ɹ������DD4�DDDaD�LD@@@@ @ @ ��۔D DDD@I���������d@�����ٴ���i�D4dDDDDDD@DDD@@D D D @���Di �@a����������� �����y�������4D�DDDDFD@DDDDD@ @ D ����� DD�K����������Di��������I����LDDD`@DDDDDDD@@D@@@  @@@ۑ�DKDD=�����y����O��9������I����D�N@DDddDF@DDD@ @@     ���lD@@DD������9����O��������@������LDDDDDDDDD@ND@DD    @D ۑ�DLDD����������DF���������I���DC�Dd D`DD@D�D@ D DAD @ ����F@@DK��������O�AO���������@��L�K�DDDDD D@�d@DD��@ ��LL`����ۙ���;DNO��ۛ�����@��F�DDD  @dDD DKD  ���D� D���������D����������@����I��d@@F@@ DDDD@@@K����@ M���F@@I��������` K����������D���D��DD@D @@D@DD@ ����@@ ���LD����ٛۙ4 I���ٹ������D���N���DDDDD @D@ 9A  ����D� 4�ۛ�����������������@���I���DFD@D  DDD@@@�;��  ����Dd ��۝���ۛ��������������@I�D�����D@ Dd@@@@D@I1����@ ߙ���� K�D�۝����������������I@��Ĺ���D @@D@ DDD @�ě��4�  ����DL;�D���ۛ�����������������I�K����@D@@@4@@@ @D��A����D ��9��D��Dl�۝�����������������`������D @K D@D9�iI9��  ����D�DDA���������ٹ���������@�������@ @D@DDDI���a�;���@ �����dAD�I�������ۛ������9�����D���<d@D D @ DDD�<�KD��1�� ������DDDɟ��۝�����ٹ���������L�ɑ���DDD D��KA�LIN<@ �����LLDa��۝��ۛ�����������	�������DD D @DD��DL��IdDAD ۙ�Dd��۽�����۝��������������IlDD@ D D DFDAIdLDDd��Ĵ@ ���II D���ۙٽ��������������I���I9DDD@D  F��ĴDdd�D�DDF@ K?�����DL�ۙ���1���ٹ����9K��I�����LL@  DDDIlD�F�FDD  K������D@D�۝���������ٛ�������K�������D@D @�DDldDD@DDDD D��������LK���������ۛ������i9�I��������D@ @ DDDDDDDDDD K����9ٹ�DdD�����ۑ������������9K����II<d@� D@  @DK�����{����LD�K�����������ٹ����L�I������IDD  @ DDD@@@@DdK������ٱ��DL���ٟ���������������K�K�����D D @@   @@?DdDD�����?����DI���ۙ�������������D��������DDD @  ��?��F@�����󟙙��DI�ۙ���������������ƙI������@L  @@������@�O���?;�����������������������iD�ɹ����ÜD F @ ��1?�0K�����3�������DD���������9�9���������I����9�4D@I @@@@��;���9�O����?yٱ���DD�۝���������������KI��������D@   �{�;�A��@����;��ɹDD��ۙ�������������9��IK����锔D@D@@��q��;K����Do��?�9��@N���������������KKI���ɑ�iDD@ @@9���A C���������y����DI���������9�����ÔIK���9���D@@@ ���� �KO��D��������I����������������K��ÙK�I�����iDD@ ?�� 	4�;;��[���@s������������������������I����ɖ��@@ @@�4@ �;��9����{| �������������ٙ����˜���ilDI�����D@  @ @94�����{��0;����	����ۙ������������<���陹����D@@ @D @  ;A������?��O7�9�I������9��������I���I<d����lD@  @@@ �94���?�����9���II����ۙ����������D�I���I���ˑ�Ɣ@D@     @C���9?������ ;=�9��K����������������D�ə1�I����KÔ�D D@@@ ��9;������D@	����I����ۙ���������DDA��NK������LD@@@    @@@DO�����1D     ����I��ۛ��������������NDF��I���I��@D@D A@@D@D ��D      9���D�����9������������DDNNI�����9IDD@D@@ D @@DF@ �@       ;�������ۛ�����������ɹ�KLDDI���I��l@D  @K @@@DLD@D       K��������ۙ���������Iɔ�L@@ə������D@@@@ A@ @DD       s1d DK���ۛ�������������<9DD���������D@ � @@@D@D       �;DD �����������������������������D  @ A@@@    @@  Ks�D@  ٹ�����������������IDDK�I����IL�D @�@@ @@  @@  �3F@   �������������9����L���II9��d@@ @@  @    G7�D  @	KۑI�����������9����IdC��������i�D�   @@   @  �D@  OI��陛��������9���I�ĴLI�����D�dDD@     @@@  7D @@ �I�������������I�����L������D�D@ � @@@@@@ @ w;D    @��ٙ���������������IKDD������DD@@@I@       @ ?4d @@@ O����I��������������@�����@ @ � @@ @@@@@@  �s4     	��������������ɹəKI���D�ə<������ @@	9  @    @ s�@ @ D��i��I���������Ü���DK�����@@@ � @@ @@@ @ 4@   I���I�������������Il��I�����9�D  K@  @  @  G�d  ����F�������I������Ĵ�DDK�������D 	� @@ @   �3@ @@@	���������������K�ɹK�Iᔔ�N������LD̔@  K