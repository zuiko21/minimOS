          @@@@@@@DDD�ND��@DDD@DND�D�NDDD                    @J@�����@����@NJK��������@ @@ @@                     JJJ�������DNDDA�NNN�D��D�N

JJ                    @@N KN�����@�N��KKK�@O������DDD@                    �
@@��������@N�A����DN�@���������   @                   @@@J�뻿��^�����ᴾNDK���[T��N@� NN@                   D�A��@ND����KK���ND���D���� D��                   @J@NNDNN��A���������N���N������D@�@N�@                   @@DNDDK���K�����A�KD�K���N�����                   � N�@N����NKKK����K����K����D�@�@DK@                    ��@NDO����ᴴ�������KA��K�N��ỾN@ K��                   D@NDJ@K����Nᱻ�����񴾴���D��D� D@
@N                  ��N�N����山��[�����Kൿ���� @�N@                  ���D�������������������KK��N@D@
@                    ���NDKA����K���񻵱������O��@�D �@@�@                  ��D�������������������������@@�
@@                   ���@��D�[��K�񿻿��[_�����N��A�@@@D                     ����DNK��K��[_�����������K����@ � ��                   ���� K������񻿿�񿱿���������� @ �O���                  ���JNKK���������������_��_�KK���D�D� K���                  ����@NK������������񿿱�������� D�@J@@����                  �񰻴K�����������������������[�K��@@
����                  ���O��D����������������������@D@����                  ����D������������������������� J@
@����                  ��N�������������������������� D����                  ��D����������������������������K D
 JK����                  ��K�D����������������������������D D O����                  ��D�NK�������������������������D� J O��                  �D��������������������������KNN@@@@���                  ��@��K�������������������������DD���                  �D����[��������������������������@J K���@                  ��N���������������_�������ND@� @A���                   ��D��������������������������DD D ��@                  ��K���������_����������_��@��@K���                   ��DN������������񿻻�����D�@���D@                  A��@任�������[��������������� D ᱱ��                  �ND�D�����[����[������K�����N�
@��@                  �D�N������[��������N��ᱻK@@ @����                  ��JDK�����������������K���J@�@                  �D��������[�����񱻱�KKNA��  @�D��@                   D @��A��A�������������NDDN�                    ������ự���[��ᱱ�NAKD�K� NO��                  D ��A���K��[���K���N��K���D @D��O�                   JND�����䱻��������K���ND��ND�ND�D
����                  �@�KAKN��������A���NNDDK��D�K��                  J��K�DA�������䱴��NKDKN��@�KD����                  ��@D�N ND��[A��ỻD�D�DDDD�@�@���                  �K����NNA�K�K���ND@���@�@K���                  �����KN�ᱱDND뱻K��뱾D @D�@    N�_�                  �N��@KK��K�����D���K�D  ���@D� @����                   [��K�����D�O��ự� D��D@@
@D�[���                  �K�@N������ND��� NKKJD
@@J@  K���                   �D��������D࿻���D���ND@@@��[���                  �@K�����J@DNA��D�_N@ ND�@DJN�@@@@K����                  �NN����    ��N����ND@    @D �����                  D�NKD���@@D��@@N�����@�  DJ@ @��@����                  @ND���K�� 
 �K���[@D@�
@ �@J @D����                  �DD�������D��K���� �@ �� @@�仱���                   D N�D���������K���������NDD�@@@@D�����                   ��DD� �������������[DN�����N�ND N����                   @�@DN���������_�������N�[�D��N�@�_���                  DN
 �����������������K����ᴻK�������                  
JJ@J�����������������D��������KNJ@ K����                   D@@@���������������D���_����DJ@K�����                   @�@���������������N����������N @������                   �@�JJ������ᱻ��������D���������N@@�����                   D�K ������D�K�������N�����������������                  @�������K��������NN��������D@  �����                   ��@���������������������K�������K��� ����                  N� D������������������D��������  ���                   @O��@K����������������N��������D JD����                   �O[@����������N����@�����[����
N  ����                  ����K��������������������K������KD @N��@                   N��������������K��������������� @A��                   񿿻A�����������������@������D��  � @                   ￻������������������K��K������D D@�N@�                   ��[[������[����������KD任����D�@@� @@ �                  ����KD�������N�������N@DK���N@�@�@���                  �������������D��D���D�� ��                  ��[DK��KA�ND��@K���@ @A�A���DDJ@ @ D��@                  �[�N��D�NNDK�����[D @�NA����@N� ��A�                  ����D�N�NND�N������@�N �@NNDN@��  �[�@                  �����D�D@JA���[D�N@@DDD@DND ND ��K@                  ��������D
N�����A�D��J
@����D@@���KK@                  �K������� N���ND��@D��JD ��D��@                  ��������@@�����D@D�NK��ND���KK@                  �D᱿���������K[����D ᱻND�@@�D���                  �K����[�K@����ND@��@ KK��ND� A����K                  ���῿�����������N�D@@������� JK���                   K�KK��������D@�NJ�N���D����@                  @KD������������� D@@@@ND������
@��N@                  �NN��[������[�  @�K�����ND �K���                  @�����A�����������D���N��A� � @��                  ��DK���N��������NND�ND��K�����@� �K���                  ������K����������N��N��ND�@��@                  �NDK���NK_�������񱱻��D��D@@�@@�K�D@                  ���῿���D�����[�������D��NN@ DK�K�                  �K@K����@KK�[����������D�D� D �@@���                  K�A��N�K��������A�KKKN
D
  ���                  ������@NNK[���������DDDND @D@�K���                  ��D�����DDN�������A��@��� J
@  @���                  ��K[��JND������[������@D@J@@�N���                  ��JK���KD D���������������@@�� K���                  ND�A����NDN���������N@DD @ @@�����                   �@@�����@@��K���������@D @�� �@����                   NND��@�DN����������@� D@@ [���                   @DNJ��������A���������NJ@@@@@D @�O���                  �
�K���D�����������@N�@ त J@���                   @DND������
D�N[���D@@D�
D@ J@ K���                   @�DN���@@D�ự�����D � @@ @� O���                   �D@��D���������D��DNDNDJD@D@�� @@�����                   D DDN����@@DND���D��@D�J@@�@K���                   @�@JND���������NDD�DD��@�NJ@@ �@@ ����                   ��ND䴱���� �DNDD��NN�D @D J@@���O���                   @@JD��K������@DD�NAD��D��NN@� @@ @ K���                  �DNK������NAND�DNN�D@ @@�@� N D���                   �@�䴴����ND���NDND@@�@��@JD���@�O���                   DDDKK��������NND���DND @�  D�@ �����                   �JD���䱵�����N�KNDDND@��@@DJJ @���                   DJDNKK��[��D��@@�
D @�@ठ@� J@@D����         