                                                                                                                                  ������������������������������������������������������         ��������������������������  ���������������������������        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �    �����    �������    �    �������    �����    �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    �����    �������    �    �������    �����    �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �    �����    �    �������������    �    �����    �        �    �        �    �                �    �        �        �    �        �    �                �    �        �        �    �����    �    �����  ������    �    �����    �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        ���������     � ������    �    �����      ����������         ����������    �          �    �          ���������                   �    �          �    �          �                            �    � ������    �    �����     � �����                 �    �                      �    �                     �    �                      �    � � ��                 �    �                      �    �   �                  �    �                      �    � ����                 �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �    �����    �����    �    �                            �    �    ��������������    �    �                 ������������    �    � � � � ��    �    ����������������������������     �    � � � � ��    �     �����������������                      �� � � � �                                                  � � � � ��                                                  � � � � ��                                                  �� � � � �                                                  � � � � ��                                                  � � � � ��                                                  �� � � � �                                                  � � � � ��                            �����������     �    � � � � ��    �     �����������������������������    �    �� � � � �    �    �����������������           �    �    ��������������    �    �                            �    �    ��������������    �    �  ww                  �    �                      �    �                      �    �                      �    �  pw                  �    �                      �    �                      �    �                      �    � w pww                  �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �                      �    �                            �    �    �������������    �    �                            �    �    �                �    �                   ����������    �    �                �    ���������         ���������     �    �����  ������    �     ����������        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �                          �                          �        �    �����    �������    �    �������    �����    �        �    �        �          �    �          �        �        �    �        �          �    �          �        �        �    ���     �������    �    �������    � ����    �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �        �                                  �        �        �����    �    �    �������������    �    �    ���        �       �    �    �                �    �    �           �       �    �    �                �    �    �           �����    �    �    �����  ������    �    �    ���        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �              �          �          �              �        �    ���������  ������    �    �����  ����������    �        �    �                    �    �                    �        �    �                    �    �                    �        �    �����������������    �    �����������������    �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �                                                      �        �������������������������������������������������������         ������������������������������������������������������                                                                                                                                        