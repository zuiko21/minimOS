��������������������                 ����������������������������                 ��������"""""�������""""""" 33333333333333333 �������"""""�������""""""" 33333333333333333 �������"""""""""""""""""" 333�������������333 ������"""""""""""""""""" 333�������������333 ������"""""""""""""""""" 33������"��"�����33 ������"""""""""""""""""" 33������"��"�����33 ������33333"""""""333333 3��"��������������3 ������33333"""""""333333 3��"��������������3 ������333333333333333333 3����������  ��"��3 �  ���333333333333333333 3����������  ��"��3 �  ���333333333333333333 3���������  ����3   ��333333333333333333 3���������  ����3   ��wwwww3333333    33 3������"��  ���3  ��wwwww3333333    33 3������"��  ���3  ��wwwwwwwwwwww   w 3���������      ��wwwwwwwwwwww   w 3���������      ��wwwwwwwwwwww     3���"�����  ��wwwwwwwwwwww     3���"�����  ��UUUUUwwwwwwwU    3�������"  �UUUUUwwwwwwwU    3�������"  �UUUUUUUUUUUUUU   3�"������ � �  �UUUUUUUUUUUUUU   3�"������ � �  �UUUUUUUUUUUUUUU    3��������       �UUUUUUUUUUUUUUU    3��������       ������UUUUUUU�����  3�����"�� ���� ������UUUUUUU�����  3�����"�� ���� ������������������� 33�"����� ��   �� ������������������� 33�"����� ��   �� ������������������� 333�������         �������������������� 333�������         ����������������   3333333333  �����������������   3333333333  �������������������                      ��������������������                      ��������������������   �  �����  �  ���������������������   �  �����  �  ������������������    ��   �������   ��  �������������������    ��   �������   ��  ��������������������������������������������������������������������������������������������������������������������                 ����������������������������                 ��������"""""�������""""""" 33333333333333333 �������"""""�������""""""" 33333333333333333 �������"""""""""""""""""" 333�������������333 ������"""""""""""""""""" 333�������������333 ������"""""""""""""""""" 33������"��"�����33 ������"""""""""""""""""" 33������"��"�����33 ������33333"""""""333333 3��"��������������3 ������33333"""""""333333 3��"��������������3 ������333333333333333333 3�����������  �"��3 ��  ��333333333333333333 3�����������  �"��3 ��  ��333333333333333333 3����������  ���3 �  �333333333333333333 3����������  ���3 �  �wwwww3333333wwwwww 3������"���  ��3   �wwwww3333333wwwwww 3������"���  ��3   �wwwwwwwwwwwww  www 3����������      �wwwwwwwwwwwww  www 3����������      �wwwwwwwwwwww  ww 3���"������  �wwwwwwwwwwww  ww 3���"������  �UUUUUwwwwwww     3�������"�  UUUUUwwwwwww     3�������"�  UUUUUUUUUUUUU  3�"������� � �  UUUUUUUUUUUUU  3�"������� � �  UUUUUUUUUUUUUU   3���������       UUUUUUUUUUUUUU   3���������       �����UUUUUUU����   3�����"��� ���� �����UUUUUUU����   3�����"��� ���� ������������������ 33�"������ ��   �� ������������������ 33�"������ ��   �� ������������������ 333��������         ������������������� 333��������         ����������������  33333333333  �����������������  33333333333  �������������������                       ��������������������                       ��������������������  �  ������  �  ���������������������  �  ������  �  ������������������   ���   �������   ��   ������������������   ���   �������   ��   ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������"""""""���������                 ������������"""""""���������                 ��������""""""""""""""""""" 33333333333333333 �������""""""""""""""""""" 33333333333333333 �������"""""""""""""""""" 333�������������333 ������"""""""""""""""""" 333�������������333 ������""""3333333""""""" 33������"��"�����33 ������""""3333333""""""" 33������"��"�����33 ������333333333333333333 3��"��������������3 ������333333333333333333 3��"��������������3 ������333333333333333333 3�����������  �"��3 ��  ��333333333333333333 3�����������  �"��3 ��  ��3333wwwwwww3333333 3����������  ���3 �  �3333wwwwwww3333333 3����������  ���3 �  �wwwwwwwwwwwwwwwwww 3������"���  ��3   �wwwwwwwwwwwwwwwwww 3������"���  ��3   �wwwwwwwwwwwwwwwwww 3����������      �wwwwwwwwwwwwwwwwww 3����������      �wwwwUUUUUUUwwwwwww 3���"������  �wwwwUUUUUUUwwwwwww 3���"������  �UUUUUUUUUUUUUUUUU  3�������"�  UUUUUUUUUUUUUUUUU  3�������"�  UUUUUUUUUUUUUU     3�"������� � �  UUUUUUUUUUUUUU     3�"������� � �  UUUU�������U   3���������       UUUU�������U   3���������       ������������    3�����"��� ���� ������������    3�����"��� ���� �������������    � 33�"������ ��   �� �������������    � 33�"������ ��   �� ��������������� 333��������         ���������������� 333��������         �������������������  33333333333  ��������������������  33333333333  ��������������������                       ���������������������                       ������������������  �  ������  �  ������������������  �  ������  �  ���������������������   ���   �������   ��   ���������������������   ���   �������   ��   �������������������������������������������������������������������������������������������������"""""""���������                 ������������"""""""���������                 ��������""""""""""""""""""" 33333333333333333 �������""""""""""""""""""" 33333333333333333 �������"""""""""""""""""" 333�������������333 ������"""""""""""""""""" 333�������������333 ������""""3333333""""""" 33������"��"�����33 ������""""3333333""""""" 33������"��"�����33 ������333333333333333333 3��"��������������3 ������333333333333333333 3��"��������������3 ������333333333333333333 3�����������  �"��3 ��  ��333333333333333333 3�����������  �"��3 ��  ��3333wwwwwww3333333 3����������  ���3 �  �3333wwwwwww3333333 3����������  ���3 �  �wwwwwwwwwwwwwwwwww 3������"���  ��3   �wwwwwwwwwwwwwwwwww 3������"���  ��3   �wwwwwwwwwwwwwwwwww 3����������      �wwwwwwwwwwwwwwwwww 3����������      �wwwwUUUUUUUwwwwwww 3���"������  �wwwwUUUUUUUwwwwwww 3���"������  �UUUUUUUUUUUUUUUU   3�������"�  UUUUUUUUUUUUUUUU   3�������"�  UUUUUUUUUUUUUU   3�"������� � �  UUUUUUUUUUUUUU   3�"������� � �  UUUU�������UU  3���������       UUUU�������UU  3���������       ������������     3�����"��� ���� ������������     3�����"��� ���� ������������  �� 33�"������ ��   �� ������������  �� 33�"������ ��   �� ����������  ��� 333��������         �����������  ��� 333��������         �������������������  33333333333  ��������������������  33333333333  �������������������                       ��������������������                       �����������������  �  ������  �  ������������������  �  ������  �  ���������������������   ���   �������   ��   ���������������������   ���   �������   ��   ��������������������������������������������������������������������������������������������������"""""""���������                 ������������"""""""���������                 ��������""""""""""""""""""" 33333333333333333 �������""""""""""""""""""" 33333333333333333 �������"""""""""""""""""" 333�������������333 ������"""""""""""""""""" 333�������������333 ������""""3333333""""""" 33������"��"�����33 ������""""3333333""""""" 33������"��"�����33 ������333333333333333333 3��"��������������3 ������333333333333333333 3��"��������������3 ������333333333333333333 3����������  ��"��3 �  ���333333333333333333 3����������  ��"��3 �  ���3333wwwwwww3333333 3���������  ����3   ��3333wwwwwww3333333 3���������  ����3   ��wwwwwwwwwwwwwwwwww 3������"��  ���3  ��wwwwwwwwwwwwwwwwww 3������"��  ���3  ��wwwwwwwwwwww    ww 3���������      ��wwwwwwwwwwww    ww 3���������      ��wwwwUUUUUUU     3���"�����  ��wwwwUUUUUUU     3���"�����  ��UUUUUUUUUUU    3�������"  �UUUUUUUUUUU    3�������"  �UUUUUUUUUUUUU     3�"������ � �  �UUUUUUUUUUUUU     3�"������ � �  �UUUU�������UUUUU   3��������       �UUUU�������UUUUU   3��������       ������������������� 3�����"�� ���� ������������������� 3�����"�� ���� ������������������� 33�"����� ��   �� ������������������� 33�"����� ��   �� ���������������  333�������         ����������������  333�������         ������������������    3333333333  �������������������    3333333333  ������������������                       �������������������                       ����������������  �  ������  �  ������������������  �  ������  �  ���������������������   ���   �������   ��   ���������������������   ���   �������   ��   ������������������������������������������������������������������������������������������������"""""�������""""""""                 ��������"""""�������""""""""                 ��������""""""""""""""""""" 33333333333333333 �������""""""""""""""""""" 33333333333333333 �������"""""""""""""""""" 333�������������333 ������"""""""""""""""""" 333�������������333 ������33333"""""""333333 33������"��"�����33 ������33333"""""""333333 33������"��"�����33 ������333333333333333333 3��"�������  �����3 �  ���333333333333333333 3��"�������  �����3 �  ���333333333333333333 3���������  �"��3   ��333333333333333333 3���������  �"��3   ��wwwww3333333wwwwww 3���������  ���3  ��wwwww3333333wwwwww 3���������  ���3  ��wwwwwwwwwwwww  www 3������"��      ��wwwwwwwwwwwww  www 3������"��      ��wwwwwwwwwwww  ww 3���������  ��wwwwwwwwwwww  ww 3���������  ��UUUUUwwwwwww     3���"����  �UUUUUwwwwwww     3���"����  �UUUUUUUUUUUUU  3�������" � �  �UUUUUUUUUUUUU  3�������" � �  �UUUUUUUUUUUUUU   3�"������       �UUUUUUUUUUUUUU   3�"������       ������UUUUUUU����   3�������� ���� ������UUUUUUU����   3�������� ���� ������������������� 3�����"�� ��   �� ������������������� 3�����"�� ��   �� ������������������� 33�"������         �������������������� 33�"������         ����������������  333��������  �����������������  333��������  �������������������   33333333333          ��������������������   33333333333          �������������������                    ���������������������                    ������������������  �  ������  �  ������������������  �  ������  �  ���������������������   ��   �������   ���   ���������������������   ��   �������   ���   ������