             K�;���;���;�����;���������;��;�;��;;��                          ;��;��������9�9999��9���������                          K�;��;;;;;�����;�������;���;����3�                          K9�������������;�����ӱ;;��0                          ��9=3���3�3������9�;����;;�����;;�                          C�;���;99�9�99999�9���3ӛ��������                          ;�������;᳻���9������;������9k��                          K���99�;������99;�9?�������9c�                          ;���;��;>1���F3�k��;;��������4                          K;��1�������9��i;��lD�9��91��;;9��>�                          C�9y���������3�����F����K�����>��                          ���999>9��K����l><aF�99;�����>0                          K;�;�9>�ka���������δ�df����K;���                          �9��99�������;9�9;��il��d��;������                          K9����;c�<;Ö���<d�<nNK��9;���>�                          K>;����9᳴�Ilk3û���ld�dƖ��k;9;90                          ����9�;��n��k;4�NN�al�3��;��                          K9>1�������ld��44���<�N�<�d;��;�<��4                          A������9�;F�Nd���K4�kKN���L>��9�;��                          K�;�;���lD�F����6ĳ�;;;�������9�                          9㛳ô��FDlF��L<;9��;�������9;;����                          K��3�ᴳ�1�F�Dd�����l;��������;��                          K93��k�FF�ll<iki>K;����������>k�                          ��;9���dLhFF�Ö���;������������ᱱ�                          K��Ó99k��FDl��㻿��;���������k�k��                          <>;�k㓶L,ld���������������?�<9���                          A���3���FD�L493�������{���������Kn4                          ;���<<��lld�K�K�����������������<<���                          K�>;ó;NDBLLi3����������������I��<>                          ;�����4��fN;�k;��������������;6Ƽ���                          C���91���ND��3��[��������������i9c��                          ���ldNldf����������������N>9�ð                          K���3���N@FN�;3����������������KKD                          ���9��<d���d��?��������������ki;���                          9k�;<��FD�?�������?�������9����                          C�in����>F���L;�����������������i<>d                          K��i9����Ll3�������91K����3L96����                          4<;����;��dFķ�������a�9��������ᴖ�                          �Ki;�ᴟ���䳻���������;����i;;<;kid                          Id���d����i���������d����d��<n��                          >Iki�ᴻ�����?������9@�ÿ���@�l1��90                          KcÖ;<>;?���{��������Ki�����k��<<n�                          C�������9��;������������������������d                          ô���>K����9?���������;����?��ô���                          <kK<<ikK�;���������{�������?�>K>0                          I㖴�ᴴ��O�����������?�������K<6�i�                          9iN;Kd����;??�������������������4��                          ��㱳�;�����������������������9ial�0                          NiN<k��;����������?�������󶖞K�                          9>������������������������4a�d0                          IkN99<<�������K�����������������˾�                          �����<<;�?��������?��������<3Da�0                          N9������Ŀ��������?��������C�;�<�                          N4��Ƴ�><6CDo�?������{��������{�6�<c�                          �>l;kKC�<��D���������?���?���9Ü0                          a䶓d��䴴n?>������������{������c�<c�                          F�Kl�IakKKÿ������������������3�ic�D                          id�if���9��{����������?������4��                          D��A��f�FF�������������������Kc�i�d                          kDi>d�i4inK���?����������{?���4�6�K�                          C��KLKN�Ɩ�o���������1����;�Ɣ��i6                          l�N4ikKl������������><;��ln����                          �la�ᶔ�D��;�{�������?����?����L<40                          CƖ>Fl69���������������{y���d�A�FN�                          ill<��k�y�������������{yC�D�Li�0                          	a��anC�`i���?��?�������{����N�N�K�                          �AKN���C������?�����������a�F����d                          N>�4�kFl`�;�������������?�?�D�F�FN�                          ���>C�FK��������������;�tnC�A�d4��                          KncNC�NH����{���������?�D�N�d�䱴                          �A���>@F����?;����?;�@�@dNCFN0                          C��>4�d$�����k����9;{���<F�F�F��@                          KFôF@��d`�����D���96��1��@hF�Dd�Di�                          F��d�dD$��?�?��@i;;��l��@�$��D�d`                          ��f�d���`����>C�;;C��@$ `�@`BFFƐ                          �d��`@`Ć�����lc�����LlF��F$�d`                          D$`@D$D$d��C������4���@`BB@F$�fƐ                          J@�d���N@?�@K?���?�C��`d`$@d�l0                          $�B@N��O�o��������B�d �,��ND�                          �JD`BDD��?�����k��@@JF�B@d$D$N`                          �@H,�@F滓������4H@HDL,D�                          FB��$$`L$���??�����HBBF@`F�F�                          �d�d$@@�Ą`@`K������?���$$�h@@$�D�@                          @d�@(BBBF�h@K�����������@B�$�@�Fd�                          �$�,$B$`ÿ����������`� �$�HF@                          D�D@@l$�LD���4������DhF@d$`                          @��@h`@@d`nFĻ������C����FH@�@�B�                          FD�D��D BC��@����������  @B�@                          �Ƥ$@�`@B�FD�N� �?������`�BJB�JB@                          `d@�D$�` B�BN��?��?����`� d�                          LB�L�@�Dl`FN`DO�������{�`dFH�B@                          $$D d`B��d�H �����{��D �h@$D �@                          �ĠDh@d�$Hd@���{�����hd$��hd$�                          BBF� FĄ`��@JF`����{��K�� @d D @@                          d�L@``FJN@dN��{?���A�l N @�                           Fd $�L��`N,$@??�����K���@d� @@                           ��D�@BFD�D$D$N	������d���HN @@F��                           `d$�$,D�H`F�$BD���������$�,@                          ��@@@�@$F�`hNF�@������?��`@K@�``                          $�@JJBD,D�F$ D$)�����{���B�DF ��                           $�@hd�BF�`���F��������F i $                           �@�$�@D@��@Dd���?��{���d�D@                          $@JD�JB��B@d��O��������d�LB�@J@                          @� d``�$�BNK��?�����`��,$@                          �HHd,@@`L`F�d$�������D � H`                          @@@`d�@d,`N `� k� Fó���9`��D�                          D
@,lJF�@N@BDl@d�D @D�`� � ``                          Dd@F�D@�@LNB@��Nd�Fn`Dd@                          @BJBJD�d�$�$, LBDd��;��HiBD�`                           `,`F�BD`�FFFF���??���� �FH@                          D@�`d@N����@Ƅ��d�K����`� Ld`                          (@��`Hd d@`�`BFF@�O����F@k F@d@�                          @(l`D@�`JBF��B�d,@D)?�0@����Hl`                           D(@@�
FDl$JD �BF@l`@N�?��`� @@D@                          �@@d,D,LL,lLd,`�d�L$D�`���d�                          DFJ@``FJBBD�F�f�D�B@�F`d��@                          �FdND�HDLlhf�FHD�@��D��FND���`                          @D��d�D�DdndFFDld�FdNDFD$DN�n@��D�                          F�F�D�D���NLlNF�llNFNl��n�F�lBBD`�@                          lD������lNF����ld�D����do�ND�klNND�             