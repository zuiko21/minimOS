""""""""""""""""""""""""""""""""""""""""""""""""&&&"b&"bb&b"b&b&""""""""""""""""""""""""""""""""""""""""""""""""&f&&"b"bb&&&&&&&""""""""""""�"""""""""""""""""""""""""""""""""""&f&"b&"bb&&&f&&"""��"""""""""/"""""��"/�""""""""""""""""""""""""&f&&"b"fb&b&&&b&"/"��/��/"//�/""��/""���"""""""""""""""""""""""""""""""""""""""""///�""�/"/"�///"/"""�"�"""""""""""""""""""""""""""""""""""""""""//��"/"/"/"�/�/"/"��""�"""""""""""""""""""""""""""""""""""""""""/""""�"/"/"�/�/"//""""�""""""""""""""""""""""""""""""""""""""""""��"/��"��/�//"��/������"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""���""""""""""""""""""""""""""""""""""""""���""""""""""""""""""",�����""""""""""""""""""""""""""""""""",�̈���""""""""""""""""""Ȉx������""""""""""""""""""""""""""",��Ȉ���x�""""""""""""""""""ȇw��������"""""""""""""""""""""""��Ȉ������s�""""""""""""""""",��3x����������"""""""""""""""""��̈�����sh��3��"""""""""""""""",�s37x�����������"""""""""""",�̈���f���w6(��38�""""""""""""""""ȇ333w���w6���������"""""",��Ȉ����f6���sb��s38�""""""""""""""",��36ffh��wwh���b������""��Ȉ����ch�wr���sb��s36��"""""""""""""",�s36b����33x���3b������̈���h���w(�g2���v(��s3f��""""""""""""""ȇ33fb���76cv���7s(��f����f�7h���s(�g2���v(��33f(�""""""""""""""ȇ36f(���sff7���76(��g6��cv�s(���s(�g2���v(��36f(�""""""""""""",�s3fb����sh�gh��76(��gr��72�s(���s(�gs���v(��3fb���""""""""""""ȇ33f(����6h�cx��76(��g2��g2�s(���s(�g78��v(�s3f(���""""""""""""ȇ36b����76h�fv��76(��g2��g2�s(���s(�g38��v(�s6f(���""""""""""",�s3fb����sf��f3��76(��g2��g2�sh���s(�g3x��v(�36b�����"""""""""",�36f(����sf��&ch�76(��g2��g2�w8���s(�g33��v(�33(�����""""""""""��36b�����6,���c<�76,��g2��g2�sv��g3,�g67��v,�c3,�����""""""""",�s3f)����76)���c6�76)��g2��g2�sv��g3)�g2c9�v)�&39������""""""""-�36b�����76)���c2�76)��g2��g2�ss��73)�g2cy�v)��c7������""""""""��36-�����72����c2�76-��g2��g2�s7m�s3-�g2f=�v-��&3}�����""""""""��33������72����c2�76-��c2��c2�37m�s3-�c2&3cv-���c7�����""""""""-�37�������r)���cb�76)��c2��c2�3g9�v3)�c2&c3v)���&3w����"""""""",�c3y������s)���3)�76)��c2��c2�3&y��s)�c2"c3v)����c7y���"""""""""�c37������72���6,�76,��c2��c2�3&s7�s,�c2�f7v,����&3w��"""""""""",�37x�����cr���2(�76(��c2��c2�3&gv�s(�c2�&7v(����s3f(�"""""""""",�33w�����cs(�gb(�76(��c2��c2�3(gv�s(�c2�&gv(����33f(�"""""""""""�c37������7(�s"��76(�h&3��3b�3(c6�s(�c2��cv(����36b�""""""""""""Ȇ33x�����72#v"��76&7(�g8�v(�3(c6�s(�c2��fv(���s36(�"""""""""""",�337�����cr'2(��737s(�f7sf(�3(&b�s(�c2��&6(���33f(�"""""""""""""�c37x����cs7b(��77s3(�"ff"��3(&b�sf�c2��&6(��s33b�""""""""""""""�c33w�����7s"���33ff(��""���f(�h�swhc2���6(��336(�"""""""""""""",�337x����36"���6ff"(���̈��"��(�ff(c2���f(�s33f(�"""""""""""""",�c33ww6��c6(���b"�����""��Ȉ����""(c2���&(�s33b��"""""""""""""""�c337sh���f���������"""""",��Ȉ���("b������336b�"""""""""""""""",�336h�����������"""""""""""",�̈���"�����s33f(�"""""""""""""""",�c3h����������"""""""""""""""""��̈������336f(�"""""""""""""""""�c6��������"""""""""""""""""""""""��Ȉ���fc6b�""""""""""""""""""Ȇh������""""""""""""""""""""""""""",��Ȉ�ff(�"""""""""""""""""",�����""""""""""""""""""""""""""""""""",�̈�(�"""""""""""""""""""���""""""""""""""""""""""""""""""""""""""���""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""")")"""""""""""'""""""""""""+�""""""""""""""""""""""""""""""""""")")"""""""""""wr""""""""""""�""""""""""""""""""""""""""""""""""")))""""""""""'''""""""""""""�""""""""""""""""""""""""""""""""""")))"""""""""""'"""""""""""""�""""""""""""""""""""""""""""""""""""��"""""""""""'""""""""""""+�"""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""")�")�"""""""'"""""'""""""""+""+"""""""""""""""""""""""""""""""""�)")"�""""""r""""""r"""""""+""+"""""""""""""""""""""""""""""""""��")"�"""""'ww"""'ww"""""""+""+"""""""""""""""""""""""""""""""""�)")"�""""""r""""""r""""""�+""+"""""""""""""""""""""""""""""""""�)")�"""""""'"""""'"""""""+�""+�""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""��"""""""""""'""""""""""""�+""""""""""""""""""""""""""""""""""")"""""""""""""'""""""""""""��""""""""""""""""""""""""""""""""""""��""""""""""'''"""""""""""�"""""""""""""""""""""""""""""""""""""")"""""""""""wr"""""""""""��""""""""""""""""""""""""""""""""""")��"""""""""""'""""""""""""�+""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""wwwwwwwwwwww"""""""""""""""""""""""""""""""""""""""""�))))���"""w"'"rw"w"w"'""""""�"�""""""""""""""""""""""""""""""")"))))")""""rww'rw'rw'rw""""""�"�""""""""""""""""""""""""""""""""�)�))�)""""w"w"rw"rwwrw""""""���"""""""""""""""""""""""""""""""")))))")""""ww''rw'rw'rw""""""�+�""""""""""""""""""""""""""""""")�))))")""""r"w"r'"w"wrw""""""�"�"""""""""""""""""""""""""""""""""""""""""""wwwwwwwwwwww""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""wwwwwwwwwwww""""""""""""""""""""""""""""""""""""""""""")��""""""w"'"'r'r"w"'""""""�"�""""""""""""""""""""""""""""""""""""�""""""rwwrw'rrw'rw""""""�+�""""""""""""""""""""""""""""""""""")"""""""w"wrw""r"wrw""""""���"""""""""""""""""""""""""""""""""""�"""""""ww'rw'rrw'rw""""""�"�"""""""""""""""""""""""""""""""""")��""""""r"wrw'rrw'rw""""""�"�"""""""""""""""""""""""""""""""""""""""""""wwwwwwwwwwww""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""'wwr"��"'wwr""""""""""""""""""""""""""""""""""""""""""""""""""""w"'w(""�wr'w""""""""""""""""""""""""""""""""""""""""")")""��""""w'rw"""�w'rw""+"���"+��"�"""""""""""""""""""""""""""""��")")""""w"'w"("�w'rw""���+""�"���""""""""""""""""""""""""""""")"")""""""w'rw"�"�w""w""���+""+"�"�"""""""""""""""""""""""""""""��")")""""w'rw(��"w'rw""���+"""��"�"""""""""""""""""""""""""""")")""��""""w"'w"�""w'rw""���+""�"�"�"""""""""""""""""""""""""""""""""""""""'wwr"(""'wwr""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""""