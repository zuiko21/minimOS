                        D@DDD��1�;��;9���D D                                         DDD�C�i�9�?1�9����� K @                                      FDDKD�1;��3�;�{���DDD@                                    D D�9A���3A��d�O��D�@                                  @DFDK�k�419�4;49k;99?���Kd  @                              @@LD�L1��4Ó;�C�c�;�D�@                                D�D�K;d1aDc��;���D�@                                dDDF���<C�DD4d;DdO��A�����4�                                D�C�K��Dk;4ddD4a3D31A;;;;a�D@                            @ @��91�d4dD4FDC@C�c@DD1���F�D                            D  �	;D�D14CDFDdd;;D0ddC���9��                           @D DC�K�91dND4Dd43D�4F�C4k�;;��D@                      D  DD�DKKDiA1�@FC���F4d44C�?���CAD @                    D DDDDDKD�DDd�DDC@31Fi;9� KK���;��� @                    @DDFF@O�D�@K` d4C�CdD1�KA6@��9@	�                    DDF�DDA@�F 4@ DD��Cc��D3F����A;O�DD                   DDdDADD@D@DDDD`c@ dc�K;�;cDF3������ D                 DKC�D`F ad4DFA` D@A4 DA�6FFF49;�����@                DDdD��d@D@ 4 D  FD	4Ad;1�d4<1dFF��;�;��9D                DdD;D@DaFD D@F� DdD4cCDDC��Fadd��{?{�4��D @            @�DD�D@1DA� @a@ cDc�DD@@c�1Ddac���������4� D           @d<da��D�Da�  F ;@D;DC6�d��1C�3����;�����KDD          DIADD4DdA`D   D4CC@<@O��a;����;91?;?������AND          @@FKALDdD4N@    @FCDa� aD adDD11C�3��3����;�{���D        @@@4FD4�d�`     ddC@4F`@DdfFF;sC1c�4�?��?���4�DDD        D�Da�C�A@    DDDD<@DAd@C dFAad4�i4�k���������K�@      @DD<4��D� @   d4C@ddD@D4F 441adC�;19;���;��;���9�     @ @FD�Dd0�@@ D` D4DFDdd@4` C�FDc�;?�=;���󱴻�    @DD DôK4F@dDFCD Ddd`dDDFDd4@@kaa�C4���;������;�d    ` dd@D���FFDDF@adFDFDDFFFDdDa @A;34a���3���?;�?�o�     @ DFDK��DDC D4�DddFF@DdCFFFDD`D�36;3�����?����@    @CdD����FFC CDF@DFDD4FF69d44dfDc���cI6k9;3��;����?�A     DDd�k�91DDDDF4FD @DdcF11���a41c��k3�6F����;�?�����     dCd1���@acA@@D@ FDd<4k63;;3���K3��;�C;4;;?��??���A     DiD;���4ddK0 D` daai1�;�������1����41�;��;3��?���I;     CAc�A�DFD16@ CD dF;3;{�����;1a��3�c3�k;1;;�����{3K     lNLd���DK�   dFFaᳶ�����{��{?3;311�3�9?4����??���i@   @AadD�K1FC   F@DdF1�{{{������3�>�3�3;���;������;    DFD4C�CA���9dd  A@dFK;;;����������3�31;4���񳳳�;3����4O�   DlL94��3�FD@  dDdD3��{����������3����;13�;��������O�   F�dCK㑳1aDD@d   Fdk3�����������7��3����11;?�������K�   K4D��4�KDad  @   DdFC3�����������1�c�;1����;�����?��  �A��O�K1CCDF@ D@ DdFDC���7��{�����󳳳3fC�93C����?����O� �Dk��D�D�CFD@ ddDFD@F3;??����������4k91K;��;�;�������@ �CCDK1�ddDDF@DDdd@ di3�������������;33�4�O�k{1���������@ `D�DaK�A�Fd DDD@F����{�������3���c;?���;�������FD  �dD4�a��iDd@  F@D ac;7?���{�������3�;A�7�?���?����ID  DDD4dAd`d  ddDdC���������������{333??�1����?������; DFC��Ka��C@d4@FD`   FDd3;??�{������?�3�����3K�11��?����O FA�K; DCFDd@D   c�������������?���3;4?����F?�3�������  �d4K�3�46FF@FDf@ @ 61;{;33;���������3�F3��3��;��??���9� 3C����DDa44F4    D41���adaa3;?���{36Dk1c��󳱳�3����@�Dad��1�dC�@aFDD`   ck>;D�FDa;{��DDF3FKf��;?������DDD��L99�KFFFD@40C`@   Ca;;���36���66f4;;1�3;?;���??����@�Dd1����I4FFD k@@  F��;�{����6?�{1���33�K���??�{����?@D��L1�9<F3ddFF� `  ac3�33333?{;;{��;�4Dd�;�C3�;3��?��?���D�DK����d;DDF@C� D  6���D@ D��;��{s1@  �{4��?��������@�DK�3�4D4f@ 90d` ;;�d   3��{��`0C�;�31���?������D�DI91�4���;44`C@C@D ak;;{��Oc�3s�3� �o;�3�o����������@DK�KCē�C��DdF�d4FF13��{>4 ��?;�?����C��k�4O�3�������?���D;91�d4FF@C1CFD@FF;{��k�;;�7��;;1��;�;���?{?�?����@��aai����iFDdd�DfFD6c�����;;3��;�{�?���?;��c���;?�������4 �;D���;CFDd6FAadcDdFD1;;�?������{�����{{���D?�1;;�����@��1��aId@DAddd4C@dcF����������3�?��{���{��F63���33����ӓ��K��A3�CDddddFFDdBFFF33�?��������{{���?���?�C��c14�����?���1񱱱�id4D@D4`dDdFDD4dF�?���{{�{?������{�6F43����;3������䔱��A4�FFFFDDfFDd FC3�{������{{{���?���?�CF3�?�;;����46������F�4dDD4$4 `   CK7�?���󷳻{��?��?16C�����������K�����1ACD4 fFF d4@@ d3;?���?���;{������{�d�df;�;�;;9;{?��CC9�;FKF@ Dd@ 6F  93������������?�{?�{CdcA��3��?�������L9�C�a�aCA@FCF`C@ d DF;3�������3�����{�??�D;�;��?����??���d�9A�4CDdKF d4dD`d0 D@dF3?������;;�������{12A;3�?���;���������K��FF4DF4@f@FFFF FFF��;��{;?����{??7�09fD;�;�1�;���1��K�9a�a4D�FC�6@DFFD`FF1a;7�������{�;���{FCd3��;{�?�������4DddDd4FDdf @AdFDdF63�?�����7�3�;??�� da4?;�?���9?����1���D1ad`aDdD FFDa�C�3{?�������3����7� N6�3�?�����������49�Da�DF@F@@@d4C1dc������?{;{�?��s�0 dd1��?�?�;������K9;9��4dF4dd`�D`BD@cFF;33;{�������{�`DFF33����?��?�?�?����K;�CDCF d@D`fC`aa��3���???���?���@FD�C?;19?;?�?�����9��6Da�Ddd�FDdd`FDC�33�3�������?{3?;{@`Dc4a;33�������󿴴�1�F�K1fDF1DfF@d4a�c��C�??�?{363�fc;�� fC�1�;������A�I944d4kA�@DdFDc0 Cc3;;s{{3ffffbfc�tFKd3;3;��?�?��;;CK�a��@C�fDc�fBDBFDFc����f&fffcc3���ddk4��3�������;�d@Ca��4FFK@@dadFF0ddc3;3�{66333����?0Daa�����?�;������;9i����F�dda30ddf;dCFFC1���;{�������3;{�@daa;{3���{3����{��DKa�;Da;DFCD4dCCdF44d4cC33;7�;33;;33��� $FCF3��?�;?����;�FC����CDC2CC�@Fdd4CFFF;;3�s��333c���� DdkF��;��;s��������D�9�I;1�;FK�dK4�BCFCfDfFacC61���;�;;{?�?� $dAa63���?����FC�C��K�CC�3CDF1dDddacFF>;;{7���������` dfF�;�;�a1k{�?�1���D�D��414aD;D�D6A�4dFF344333��{{�?��F FDc3�3����������A4dA9;�D`C3a�6Dd;�3Fd4aicfF;;s��{�����dBD K�4?�3��?���;��FFDaKFDCFD3�D34C@�C�FF61acc33�?������?0FDdFDCvF?3;����;���� DCNDd;Fddi4c��4d33F4FFc�661a;;3������{�ddFF�1�K13;�����9�� 3�D44FC1FF4dFd1�FD4afFFC3Dk;663���7�����DFD`dd��;3��3����;;;F ��;6ddDF496CdcDd3d3DF46K63;133;3�?;;�`BFFFFC3���;;�???����<4K3�IFDDCFA�4Fc�cF6CddfC33C3��;;3�;3��0dddFDdk;;7�;?;�?�����6ca6F4DfCFD6�3A3Ddac�63��3�3;3�3FD d4FDd`aa�;�C�������O�I;�D<1DFFd9cCcC3FfC6;1k�C;;�;�3�;4CFFddddFFF�;;3��?����;OD�13CfFDdCDd�c�3dCcC��;;3�;�s�3�da�d`CFDdd43�;;?�;�������O�C�A��Ddda3;;3444666C33�3;3�3��3�FFDdddFFFF3��;��;�����9O��I�1�1aFfDf�334;6F1;���;󳳿s�?;��FCFFF4d44ak13��������?�d��F�㓓�4DdDd4��364f�;;;;3;3�{;w��Di4add4CFC4���������@�0A�kaddFcFd3�3;3�3c;3?6c�3�??��?3dF�FDdDd4c��;;;;?����9�@K�FAf�A4dFc;;3;3����;�1;?�3󷷳�{;CKd94FDfCa�3��3�??�����1`C��46F@f36�33;3;3��3�3�333�?�;3���;�F��dfd4;����������L@Daa�a�d93;;;;;3�;4;3;34;{;���;{{;;K4a4CAc6a3;;?;43��{�����0 DC<3;3�����;33�;;;;c3��3���;91�9id�<adi969����������91� FC�da�33�;;??;7���?����{�33�3?���C3�CKCCCF31�3�;;4a3����;�K`@D�FD;4��;������{{3;�?��?�3��;����DKCFFF44c�3��;�;3����DD@9Ca��33;3;???;�����;�����s�s3���FD94d4dcCFa;�3;C�;?�N@4d3K3c��;���������;?����{�{�?��33316FCKFDd4C3�;;�c���O��  FD�K99;3�3�?����?;�;�;{������?�����D4a�c3fc�3��;913�4O�4  A�dC4�33���{���������?�{?�����337�;;49c�;�3��񳳔�ƳO0 �D��;;�;;;��������7�k�{?���?���?;1�dCcK3i3�C�?;;3;C��� �4A�c3;;{?�������?;6�{�����?����;;{>�d��c�?4;;��C��3C��`4@�4��������������������s�����?���{?;a�13CcC����D09dd�  ` �c3;;{?�����������{�7�{?;;?�������󳓳;4k�Da?�3����@�K0   F ����;?;s��������?{�?�{{;{{�������?3C��1F6;����9@4CdD   `O�c;3����?��������?�;���??�������3��4D�7�?�;K4  K    @�C�;;?{���������{{����{�����������;34;;�C6;��3��;@  �6D    �;;;;{{���������������???;���������C���KD�33���B   �>@   �333����{?�����?{K�C�������������;6��4c3K3�;0B �dd  O�i;;;{{{?���������������{������������3;��C�a13;9�D@   FD  �c33��;{����������?{����7�7���?������3��d;;��K��$  ` F  ���;;�{{�����������{o�;��{��{;�������;;;�CC�c�3�O�D        ��3;3���;����������{{�4����������?�����;6�F93C��K�0        �6��??;{{{?{{{����{������?;?�����������;3�3�;��;;;3��       ���33����������?�??���k3�������?�������3�?�43�;A�D`      